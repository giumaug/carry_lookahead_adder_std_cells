magic
tech sky130A
magscale 1 2
timestamp 1695892320
<< nwell >>
rect 566 269 597 590
rect 1213 269 1238 590
rect 650 -399 704 -78
<< locali >>
rect 537 535 564 569
rect 600 535 634 569
rect 1172 535 1210 569
rect 1245 535 1271 569
rect -10 135 50 150
rect -10 100 10 135
rect 44 100 50 135
rect -10 90 50 100
rect 527 -9 565 25
rect 600 -9 634 25
rect 1173 -9 1210 25
rect 1245 -9 1272 25
rect 624 -133 660 -99
rect 695 -133 734 -99
rect 560 -350 570 -310
rect 757 -371 791 -337
rect 622 -677 664 -643
rect 700 -677 733 -643
<< viali >>
rect 564 535 600 569
rect 1210 535 1245 569
rect 658 296 694 330
rect 212 223 246 257
rect 340 223 374 257
rect 468 223 502 257
rect 852 223 886 257
rect 980 223 1014 257
rect 1108 223 1142 257
rect 1492 223 1526 257
rect 1620 223 1654 257
rect 1748 223 1782 257
rect 10 100 44 135
rect 565 -9 600 25
rect 1210 -9 1245 25
rect 660 -133 695 -99
rect 572 -355 606 -320
rect 19 -445 53 -411
rect 165 -445 199 -411
rect 280 -445 316 -410
rect 380 -445 415 -411
rect 760 -470 795 -435
rect 951 -445 986 -411
rect 1080 -445 1114 -411
rect 1208 -445 1242 -411
rect 664 -677 700 -643
<< metal1 >>
rect -150 585 -7 600
rect -150 530 -135 585
rect -80 530 -7 585
rect -150 504 -7 530
rect 534 569 635 600
rect 534 535 564 569
rect 600 535 635 569
rect 534 504 635 535
rect 1175 569 1273 600
rect 1175 535 1210 569
rect 1245 535 1273 569
rect 1175 504 1273 535
rect 1803 504 1860 600
rect 640 330 710 340
rect 640 296 658 330
rect 694 300 1660 330
rect 694 296 710 300
rect 640 290 710 296
rect 450 270 540 280
rect 195 257 260 270
rect 195 223 212 257
rect 246 223 260 257
rect 195 204 260 223
rect 320 257 390 270
rect 320 223 340 257
rect 374 223 390 257
rect 320 200 390 223
rect 450 200 460 270
rect 530 200 540 270
rect 834 257 900 270
rect 834 223 852 257
rect 886 223 900 257
rect 834 204 900 223
rect 970 257 1020 270
rect 970 223 980 257
rect 1014 223 1020 257
rect 450 190 540 200
rect 970 150 1020 223
rect 1090 260 1170 270
rect 1090 200 1100 260
rect 1160 200 1170 260
rect 1475 257 1535 270
rect 1475 223 1492 257
rect 1526 223 1535 257
rect 1475 210 1535 223
rect 1610 257 1660 300
rect 1610 223 1620 257
rect 1654 223 1660 257
rect 1610 211 1660 223
rect 1740 260 1820 270
rect 1740 257 1750 260
rect 1740 223 1748 257
rect 1090 190 1170 200
rect 1740 200 1750 223
rect 1810 200 1820 260
rect 1740 190 1820 200
rect -10 135 1020 150
rect -10 100 10 135
rect 44 120 1020 135
rect 44 100 59 120
rect -10 90 59 100
rect 533 25 634 56
rect 533 -9 565 25
rect 600 -9 634 25
rect 533 -40 634 -9
rect 1176 25 1272 56
rect 1176 -9 1210 25
rect 1245 -9 1272 25
rect 1176 -40 1272 -9
rect 1818 40 1960 56
rect 1818 -15 1880 40
rect 1935 -15 1960 40
rect 1818 -40 1960 -15
rect -150 -90 -7 -68
rect -150 -95 0 -90
rect -150 -150 -135 -95
rect -80 -150 0 -95
rect -150 -155 0 -150
rect 622 -99 735 -68
rect 622 -133 660 -99
rect 695 -133 735 -99
rect -150 -164 -8 -155
rect 622 -164 735 -133
rect 560 -320 615 -310
rect 560 -350 572 -320
rect 563 -355 572 -350
rect 606 -350 1120 -320
rect 606 -355 620 -350
rect 563 -370 620 -355
rect 140 -390 230 -380
rect 5 -411 65 -395
rect 5 -445 19 -411
rect 53 -445 65 -411
rect 5 -460 65 -445
rect 140 -460 150 -390
rect 220 -460 230 -390
rect 140 -470 230 -460
rect 260 -410 330 -400
rect 260 -445 280 -410
rect 316 -445 330 -410
rect 260 -460 330 -445
rect 360 -410 440 -400
rect 260 -500 300 -460
rect 360 -470 370 -410
rect 430 -470 440 -410
rect 940 -411 1000 -390
rect 360 -480 440 -470
rect 745 -435 809 -420
rect 745 -470 760 -435
rect 795 -470 809 -435
rect 745 -495 809 -470
rect 940 -445 951 -411
rect 986 -445 1000 -411
rect 220 -510 300 -500
rect 220 -570 230 -510
rect 290 -570 300 -510
rect 940 -520 1000 -445
rect 1070 -411 1120 -350
rect 1070 -445 1080 -411
rect 1114 -445 1120 -411
rect 1070 -458 1120 -445
rect 1195 -411 1260 -395
rect 1195 -445 1208 -411
rect 1242 -445 1260 -411
rect 1195 -460 1260 -445
rect 1290 -480 1370 -470
rect 1290 -520 1300 -480
rect 940 -540 1300 -520
rect 1360 -540 1370 -480
rect 940 -550 1370 -540
rect 940 -551 1290 -550
rect 220 -580 300 -570
rect 627 -643 734 -612
rect 627 -677 664 -643
rect 700 -677 734 -643
rect 627 -708 734 -677
rect 1277 -630 1960 -612
rect 1277 -685 1880 -630
rect 1935 -685 1960 -630
rect 1277 -708 1960 -685
<< via1 >>
rect -135 530 -80 585
rect 460 257 530 270
rect 460 223 468 257
rect 468 223 502 257
rect 502 223 530 257
rect 460 200 530 223
rect 1100 257 1160 260
rect 1100 223 1108 257
rect 1108 223 1142 257
rect 1142 223 1160 257
rect 1100 200 1160 223
rect 1750 257 1810 260
rect 1750 223 1782 257
rect 1782 223 1810 257
rect 1750 200 1810 223
rect 1880 -15 1935 40
rect -135 -150 -80 -95
rect 150 -411 220 -390
rect 150 -445 165 -411
rect 165 -445 199 -411
rect 199 -445 220 -411
rect 150 -460 220 -445
rect 370 -411 430 -410
rect 370 -445 380 -411
rect 380 -445 415 -411
rect 415 -445 430 -411
rect 370 -470 430 -445
rect 230 -570 290 -510
rect 1300 -540 1360 -480
rect 1880 -685 1935 -630
<< metal2 >>
rect -150 585 -50 600
rect -150 530 -135 585
rect -80 530 -50 585
rect -150 -95 -50 530
rect 1210 350 1770 380
rect 450 270 540 280
rect 450 200 460 270
rect 530 200 540 270
rect 450 190 540 200
rect 1090 260 1170 270
rect 1090 200 1100 260
rect 1160 200 1170 260
rect 1090 190 1170 200
rect -150 -150 -135 -95
rect -80 -150 -50 -95
rect -150 -710 -50 -150
rect 460 -180 500 190
rect 160 -210 500 -180
rect 160 -211 470 -210
rect 160 -380 190 -211
rect 1100 -260 1130 190
rect 260 -290 1130 -260
rect 140 -390 230 -380
rect 140 -460 150 -390
rect 220 -460 230 -390
rect 140 -470 230 -460
rect 260 -390 300 -290
rect 989 -291 1130 -290
rect 1210 -340 1240 350
rect 1740 270 1770 350
rect 1740 260 1820 270
rect 1740 200 1750 260
rect 1810 200 1820 260
rect 1740 190 1820 200
rect 360 -370 1240 -340
rect 260 -460 299 -390
rect 360 -400 390 -370
rect 360 -410 440 -400
rect 260 -500 300 -460
rect 360 -470 370 -410
rect 430 -470 440 -410
rect 1300 -470 1340 149
rect 1860 40 1960 600
rect 1860 -15 1880 40
rect 1935 -15 1960 40
rect 360 -480 440 -470
rect 1290 -480 1370 -470
rect 220 -510 300 -500
rect 220 -570 230 -510
rect 290 -570 300 -510
rect 1290 -540 1300 -480
rect 1360 -540 1370 -480
rect 1290 -550 1370 -540
rect 220 -580 300 -570
rect 1860 -630 1960 -15
rect 1860 -685 1880 -630
rect 1935 -685 1960 -630
rect 1860 -710 1960 -685
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_0
timestamp 1691611044
transform 1 0 -12 0 1 8
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_1
timestamp 1691611044
transform 1 0 628 0 1 8
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_2
timestamp 1691611044
transform 1 0 1268 0 1 8
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_3
timestamp 1691611044
transform 1 0 728 0 1 -660
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  sky130_fd_sc_hd__and4_1_0
timestamp 1691611044
transform 1 0 -12 0 1 -660
box -38 -48 682 592
<< labels >>
flabel metal2 1130 270 1130 270 1 FreeSans 128 0 0 0 P3
port 6 n
flabel metal1 870 270 870 270 1 FreeSans 128 0 0 0 G3
port 7 n
flabel metal2 1770 270 1770 270 1 FreeSans 128 0 0 0 P4
port 8 n
flabel metal1 1510 270 1510 270 1 FreeSans 128 0 0 0 G4
port 9 n
flabel metal2 490 270 490 270 1 FreeSans 128 0 0 0 P2
port 4 n
flabel metal1 1230 -400 1230 -400 1 FreeSans 128 0 0 0 CI
port 1 n
flabel metal1 40 -410 40 -410 1 FreeSans 64 0 0 0 P1
port 2 n
flabel metal1 350 270 350 270 1 FreeSans 128 0 0 0 G1
port 3 n
flabel metal1 750 -455 750 -455 1 FreeSans 128 0 0 0 CO
port 10 n
flabel viali 230 225 230 225 1 FreeSans 128 0 0 0 G2
port 5 n
flabel metal1 s 125 555 125 555 1 FreeSans 128 0 0 0 VDD
port 11 n
flabel metal1 s 123 -658 123 -658 1 FreeSans 128 0 0 0 GND
port 12 n
flabel nwell s 124 579 124 579 1 FreeSans 64 0 0 0 VPB
port 13 n
flabel pwell s 120 -695 120 -695 1 FreeSans 64 0 0 0 VPN
port 14 n
<< end >>
