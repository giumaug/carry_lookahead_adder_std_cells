ADDER

v1 CI GND pwl 0 0ps
v2 A4 GND pwl 0 0ps
v3 B4 GND pwl 0 0ps 1000ps 0 1050ps 1.8
v4 A3 GND pwl 0 0ps
v5 B3 GND pwl 0 0ps 1000ps 0 1050ps 1.8
v6 A2 GND pwl 0 0ps
v7 B2 GND pwl 0 0ps 1000ps 0 1050ps 1.8
v8 A1 GND pwl 0 0ps 1000ps 0 1050ps 1.8
v9 B1 GND pwl 0 0ps 1000ps 0 1050ps 1.8
v10 VDD GND pwl 0 1.8

Xadder_0 A1 B1 A2 B2 A3 B3 A4 B4 A5 B5 A6 B6 A7 B7 A8 B8 A9 B9 A10 B10 A11 B11
+ A12 B12 A13 B13 A14 B14 A15 B15 A16 B16 S1 S2 S3 S4 S5 S6 S7 S8 S9 S10 S11 S12 S13
+ S14 S15 S16 CI CO

Xadder_4_0 A1 B1 A2 B2 A3 B3 A4 B4 CI S1 S2 S3 S4 CO VDD GND adder_4

.measure tran tpdr TRIG v(B1) VAL=0.1 RISE=1 TARG v(co) VAL=1.7 RISE=1
*.measure tran tpdf TRIG v(B1) VAL=1.7 FALL=1 TARG v(co) VAL=0.1 FALL=1 CROSS=LAST


.lib /opt/open_pdks/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.tran 10p 204800ps
.options method=gear
.tran 40ps 4000ps
.save all

.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X a_384_47# a_81_21# a_299_297#
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.229 ps=1.57 w=0.65 l=0.15
**devattr s=10270,288 d=3575,185
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.69 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5500,255
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.69 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.69 as=0.18 ps=1.69 w=1 l=0.15
**devattr s=5500,255 d=5600,256
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.229 pd=1.57 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=10270,288
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.229 pd=1.57 as=0.091 ps=0.93 w=0.65 l=0.15
**devattr s=3640,186 d=6890,366
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.69 as=0.18 ps=1.69 w=1 l=0.15
**devattr s=5600,256 d=10600,506
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
**devattr s=3575,185 d=3640,186
C0 VGND A1 0.0786f
C1 a_81_21# a_384_47# 0.00138f
C2 VPB B1 0.0387f
C3 a_299_297# VPWR 0.202f
C4 A2 VPB 0.0373f
C5 VGND a_384_47# 0.00366f
C6 A1 VPWR 0.0209f
C7 a_299_297# A1 0.0585f
C8 a_81_21# B1 0.148f
C9 a_81_21# A2 7.47e-19
C10 a_384_47# VPWR 4.08e-19
C11 VGND B1 0.0181f
C12 VPB X 0.0108f
C13 a_299_297# a_384_47# 1.48e-19
C14 A2 VGND 0.0495f
C15 A1 a_384_47# 0.00884f
C16 a_81_21# X 0.112f
C17 B1 VPWR 0.0196f
C18 a_299_297# B1 0.00863f
C19 A2 VPWR 0.0201f
C20 a_299_297# A2 0.0468f
C21 VGND X 0.0512f
C22 A1 B1 0.0817f
C23 A2 A1 0.0921f
C24 a_81_21# VPB 0.0593f
C25 X VPWR 0.0847f
C26 VGND VPB 0.00713f
C27 a_81_21# VGND 0.173f
C28 VPB VPWR 0.068f
C29 a_299_297# VPB 0.0111f
C30 A1 VPB 0.0264f
C31 a_81_21# VPWR 0.146f
C32 a_81_21# a_299_297# 0.0821f
C33 a_81_21# A1 0.0568f
C34 VGND VPWR 0.0579f
C35 X B1 3.04e-20
C36 a_299_297# VGND 0.00772f
C37 VGND VNB 0.364f
C38 VPWR VNB 0.286f
C39 X VNB 0.0945f
C40 A2 VNB 0.144f
C41 A1 VNB 0.0996f
C42 B1 VNB 0.109f
C43 VPB VNB 0.605f
C44 a_299_297# VNB 0.0348f
C45 a_81_21# VNB 0.147f
.ends

.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X a_109_47# a_197_47# a_303_47#
+ a_27_47#
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.139 ps=0.987 w=0.42 l=0.15
**devattr s=3108,158 d=2352,140
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=3192,160
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.332 ps=2.35 w=1 l=0.15
**devattr s=12498,336 d=10400,504
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2772,150
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.139 ps=0.987 w=0.42 l=0.15
**devattr s=4368,272 d=2940,154
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.139 pd=0.987 as=0.0662 ps=0.735 w=0.42 l=0.15
**devattr s=2352,140 d=12498,336
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.154 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=7851,266
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.139 pd=0.987 as=0.0662 ps=0.735 w=0.42 l=0.15
**devattr s=2940,154 d=3108,158
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.238 ps=1.62 w=0.65 l=0.15
**devattr s=7851,266 d=6760,364
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2436,142
C0 VGND a_197_47# 0.00387f
C1 VPB VPWR 0.077f
C2 VGND VPWR 0.0662f
C3 C B 0.161f
C4 A B 0.0839f
C5 D X 0.00746f
C6 a_27_47# a_109_47# 0.00578f
C7 a_303_47# a_27_47# 0.00119f
C8 VPB B 0.0643f
C9 VGND B 0.0453f
C10 X VPWR 0.0945f
C11 D VPWR 0.0207f
C12 C a_109_47# 1.72e-20
C13 a_303_47# C 0.00527f
C14 a_197_47# VPWR 5.24e-19
C15 VGND a_109_47# 0.00223f
C16 VGND a_303_47# 0.00381f
C17 a_197_47# B 0.00623f
C18 B VPWR 0.0231f
C19 D a_303_47# 0.00119f
C20 VPWR a_109_47# 4.66e-19
C21 C a_27_47# 0.0516f
C22 A a_27_47# 0.153f
C23 a_303_47# VPWR 4.83e-19
C24 B a_109_47# 0.00153f
C25 VPB a_27_47# 0.082f
C26 VGND a_27_47# 0.132f
C27 VPB C 0.0609f
C28 A VPB 0.0907f
C29 VGND C 0.0408f
C30 VGND A 0.0151f
C31 X a_27_47# 0.0754f
C32 D a_27_47# 0.107f
C33 VGND VPB 0.00852f
C34 a_197_47# a_27_47# 0.00167f
C35 a_27_47# VPWR 0.326f
C36 D C 0.18f
C37 C a_197_47# 0.00123f
C38 X VPB 0.0111f
C39 VGND X 0.0903f
C40 C VPWR 0.021f
C41 A VPWR 0.044f
C42 a_27_47# B 0.13f
C43 D VPB 0.0782f
C44 VGND D 0.0898f
C45 VGND VNB 0.393f
C46 X VNB 0.0933f
C47 VPWR VNB 0.335f
C48 D VNB 0.13f
C49 C VNB 0.11f
C50 B VNB 0.112f
C51 A VNB 0.221f
C52 VPB VNB 0.693f
C53 a_27_47# VNB 0.175f
.ends

.subckt adder_2 CI P1 G1 P2 G2 P3 G3 P4 G4 CO sky130_fd_sc_hd__a21o_1_0/a_81_21# sky130_fd_sc_hd__and4_1_0/a_27_47#
+ sky130_fd_sc_hd__a21o_1_0/a_384_47# sky130_fd_sc_hd__a21o_1_1/X sky130_fd_sc_hd__a21o_1_0/a_299_297#
+ sky130_fd_sc_hd__a21o_1_1/a_81_21# VPB sky130_fd_sc_hd__a21o_1_1/a_299_297# sky130_fd_sc_hd__a21o_1_1/a_384_47#
+ sky130_fd_sc_hd__a21o_1_2/a_299_297# sky130_fd_sc_hd__and4_1_0/a_109_47# sky130_fd_sc_hd__a21o_1_2/X
+ sky130_fd_sc_hd__a21o_1_0/X sky130_fd_sc_hd__and4_1_0/X sky130_fd_sc_hd__a21o_1_3/a_299_297#
+ sky130_fd_sc_hd__a21o_1_2/a_81_21# VNB sky130_fd_sc_hd__and4_1_0/a_197_47# sky130_fd_sc_hd__a21o_1_2/a_384_47#
+ sky130_fd_sc_hd__and4_1_0/a_303_47# sky130_fd_sc_hd__a21o_1_3/a_81_21# sky130_fd_sc_hd__a21o_1_3/a_384_47#
Xsky130_fd_sc_hd__a21o_1_0 G1 P2 G2 VNB VNB VPB VPB sky130_fd_sc_hd__a21o_1_0/X sky130_fd_sc_hd__a21o_1_0/a_384_47#
+ sky130_fd_sc_hd__a21o_1_0/a_81_21# sky130_fd_sc_hd__a21o_1_0/a_299_297# sky130_fd_sc_hd__a21o_1
Xsky130_fd_sc_hd__a21o_1_1 sky130_fd_sc_hd__a21o_1_0/X P3 G3 VNB VNB VPB VPB sky130_fd_sc_hd__a21o_1_1/X
+ sky130_fd_sc_hd__a21o_1_1/a_384_47# sky130_fd_sc_hd__a21o_1_1/a_81_21# sky130_fd_sc_hd__a21o_1_1/a_299_297#
+ sky130_fd_sc_hd__a21o_1
Xsky130_fd_sc_hd__a21o_1_2 sky130_fd_sc_hd__a21o_1_1/X P4 G4 VNB VNB VPB VPB sky130_fd_sc_hd__a21o_1_2/X
+ sky130_fd_sc_hd__a21o_1_2/a_384_47# sky130_fd_sc_hd__a21o_1_2/a_81_21# sky130_fd_sc_hd__a21o_1_2/a_299_297#
+ sky130_fd_sc_hd__a21o_1
Xsky130_fd_sc_hd__a21o_1_3 sky130_fd_sc_hd__and4_1_0/X CI sky130_fd_sc_hd__a21o_1_2/X
+ VNB VNB VPB VPB CO sky130_fd_sc_hd__a21o_1_3/a_384_47# sky130_fd_sc_hd__a21o_1_3/a_81_21#
+ sky130_fd_sc_hd__a21o_1_3/a_299_297# sky130_fd_sc_hd__a21o_1
Xsky130_fd_sc_hd__and4_1_0 P4 P2 P3 P1 VNB VNB VPB VPB sky130_fd_sc_hd__and4_1_0/X
+ sky130_fd_sc_hd__and4_1_0/a_109_47# sky130_fd_sc_hd__and4_1_0/a_197_47# sky130_fd_sc_hd__and4_1_0/a_303_47#
+ sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__and4_1
C0 sky130_fd_sc_hd__a21o_1_2/a_81_21# sky130_fd_sc_hd__a21o_1_1/X 0.0421f
C1 VNB G1 -0.00488f
C2 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__a21o_1_1/X 0.0261f
C3 P2 sky130_fd_sc_hd__a21o_1_0/a_299_297# 0.0456f
C4 sky130_fd_sc_hd__and4_1_0/X sky130_fd_sc_hd__a21o_1_1/a_384_47# 1.46e-21
C5 G3 sky130_fd_sc_hd__a21o_1_1/X 0.0595f
C6 sky130_fd_sc_hd__and4_1_0/a_197_47# sky130_fd_sc_hd__and4_1_0/X 1.78e-19
C7 P3 G4 0.0694f
C8 sky130_fd_sc_hd__a21o_1_1/a_299_297# P2 0.0566f
C9 sky130_fd_sc_hd__a21o_1_3/a_81_21# CO 0.00936f
C10 sky130_fd_sc_hd__a21o_1_3/a_299_297# P1 2.61e-19
C11 sky130_fd_sc_hd__and4_1_0/X P4 4.68e-20
C12 VNB CO -0.00689f
C13 VPB sky130_fd_sc_hd__a21o_1_3/a_81_21# -0.0123f
C14 sky130_fd_sc_hd__a21o_1_1/a_384_47# sky130_fd_sc_hd__a21o_1_0/X 6.97e-19
C15 VNB sky130_fd_sc_hd__a21o_1_2/a_384_47# -2.27e-19
C16 sky130_fd_sc_hd__a21o_1_2/X G1 4.98e-20
C17 VPB VNB -0.275f
C18 sky130_fd_sc_hd__and4_1_0/a_197_47# sky130_fd_sc_hd__a21o_1_0/X 5.93e-21
C19 sky130_fd_sc_hd__and4_1_0/X sky130_fd_sc_hd__a21o_1_1/X 5.37e-20
C20 sky130_fd_sc_hd__a21o_1_0/a_81_21# G2 0.0401f
C21 P4 sky130_fd_sc_hd__a21o_1_0/X 5.9e-20
C22 VPB sky130_fd_sc_hd__a21o_1_2/a_81_21# -0.0132f
C23 P3 sky130_fd_sc_hd__a21o_1_3/a_81_21# 2.3e-19
C24 sky130_fd_sc_hd__a21o_1_2/X CO 0.0504f
C25 P4 sky130_fd_sc_hd__and4_1_0/a_27_47# 0.00576f
C26 P3 VNB 0.543f
C27 sky130_fd_sc_hd__a21o_1_2/X VPB 1.21f
C28 VPB G3 -6.71e-19
C29 P2 sky130_fd_sc_hd__a21o_1_2/a_299_297# 0.055f
C30 sky130_fd_sc_hd__a21o_1_0/X sky130_fd_sc_hd__a21o_1_1/X 0.121f
C31 sky130_fd_sc_hd__and4_1_0/a_197_47# P2 2.63e-19
C32 G4 VNB 8.25e-19
C33 P4 sky130_fd_sc_hd__a21o_1_1/a_81_21# 1.01e-19
C34 P4 P2 0.197f
C35 sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__a21o_1_1/X 1.67e-19
C36 P3 sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.0706f
C37 P3 sky130_fd_sc_hd__a21o_1_2/X 0.0674f
C38 P3 G3 0.0176f
C39 sky130_fd_sc_hd__a21o_1_0/X G1 0.0691f
C40 sky130_fd_sc_hd__a21o_1_1/a_81_21# sky130_fd_sc_hd__a21o_1_1/X 0.0447f
C41 sky130_fd_sc_hd__and4_1_0/X CO 0.13f
C42 G4 sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.0188f
C43 P2 sky130_fd_sc_hd__a21o_1_1/X 0.627f
C44 sky130_fd_sc_hd__and4_1_0/X sky130_fd_sc_hd__a21o_1_2/a_384_47# 1.23e-20
C45 VPB sky130_fd_sc_hd__and4_1_0/X 0.0202f
C46 sky130_fd_sc_hd__a21o_1_2/X G4 0.00776f
C47 VNB sky130_fd_sc_hd__a21o_1_3/a_81_21# -0.0199f
C48 sky130_fd_sc_hd__a21o_1_2/a_384_47# sky130_fd_sc_hd__a21o_1_0/X 1.12e-20
C49 VPB sky130_fd_sc_hd__a21o_1_0/X 0.0377f
C50 P2 G1 0.0935f
C51 sky130_fd_sc_hd__and4_1_0/a_303_47# VPB -4.83e-19
C52 P3 sky130_fd_sc_hd__and4_1_0/X 0.00586f
C53 sky130_fd_sc_hd__and4_1_0/a_27_47# CO 0.00246f
C54 VPB sky130_fd_sc_hd__and4_1_0/a_27_47# -0.0199f
C55 VNB sky130_fd_sc_hd__a21o_1_2/a_81_21# -0.0181f
C56 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__a21o_1_3/a_81_21# 0.07f
C57 G4 sky130_fd_sc_hd__and4_1_0/X 1.98e-20
C58 P4 P1 4.35e-19
C59 sky130_fd_sc_hd__a21o_1_2/X VNB 0.0224f
C60 P2 CO 4.84e-19
C61 G3 VNB 6.81e-19
C62 sky130_fd_sc_hd__a21o_1_2/a_384_47# P2 2.47e-20
C63 P3 sky130_fd_sc_hd__a21o_1_0/X 0.0694f
C64 VPB sky130_fd_sc_hd__a21o_1_1/a_81_21# -0.00647f
C65 VPB P2 0.383f
C66 P3 sky130_fd_sc_hd__and4_1_0/a_303_47# 4.7e-19
C67 VPB sky130_fd_sc_hd__a21o_1_3/a_384_47# -1.62e-19
C68 VPB CI 0.00996f
C69 sky130_fd_sc_hd__a21o_1_0/a_384_47# sky130_fd_sc_hd__a21o_1_1/X 1.32e-20
C70 G4 sky130_fd_sc_hd__a21o_1_0/X 3.47e-20
C71 P1 sky130_fd_sc_hd__a21o_1_1/X 4.83e-20
C72 P3 sky130_fd_sc_hd__and4_1_0/a_27_47# 0.0397f
C73 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.02f
C74 sky130_fd_sc_hd__a21o_1_1/X G2 1.59e-19
C75 sky130_fd_sc_hd__a21o_1_0/a_81_21# sky130_fd_sc_hd__a21o_1_1/X 0.0018f
C76 sky130_fd_sc_hd__a21o_1_2/X G3 4.15e-19
C77 sky130_fd_sc_hd__and4_1_0/X sky130_fd_sc_hd__a21o_1_3/a_81_21# 0.0697f
C78 P3 P2 0.155f
C79 VNB sky130_fd_sc_hd__and4_1_0/X 0.251f
C80 sky130_fd_sc_hd__a21o_1_0/a_384_47# G1 4.61e-19
C81 G4 P2 0.00574f
C82 G1 G2 0.0921f
C83 sky130_fd_sc_hd__a21o_1_0/a_81_21# G1 0.00416f
C84 sky130_fd_sc_hd__a21o_1_1/a_299_297# P4 1.23e-19
C85 sky130_fd_sc_hd__and4_1_0/X sky130_fd_sc_hd__a21o_1_2/a_81_21# 4.69e-20
C86 VNB sky130_fd_sc_hd__a21o_1_0/X 0.461f
C87 sky130_fd_sc_hd__a21o_1_1/X sky130_fd_sc_hd__a21o_1_0/a_299_297# 0.0315f
C88 sky130_fd_sc_hd__and4_1_0/a_303_47# VNB 3.12e-20
C89 sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__a21o_1_3/a_81_21# 0.0108f
C90 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__and4_1_0/X 0.132f
C91 sky130_fd_sc_hd__a21o_1_3/a_299_297# VPB -5.68e-32
C92 P1 CO 0.00943f
C93 VPB sky130_fd_sc_hd__a21o_1_0/a_384_47# -3.87e-19
C94 VNB sky130_fd_sc_hd__and4_1_0/a_27_47# 0.00805f
C95 VPB P1 0.00652f
C96 sky130_fd_sc_hd__a21o_1_1/a_299_297# sky130_fd_sc_hd__a21o_1_1/X 0.0338f
C97 sky130_fd_sc_hd__a21o_1_0/X sky130_fd_sc_hd__a21o_1_2/a_81_21# 1.2e-19
C98 VPB G2 0.0175f
C99 sky130_fd_sc_hd__a21o_1_3/a_81_21# P2 6.76e-19
C100 VPB sky130_fd_sc_hd__a21o_1_0/a_81_21# -0.00151f
C101 sky130_fd_sc_hd__and4_1_0/a_109_47# VPB -4.66e-19
C102 VNB sky130_fd_sc_hd__a21o_1_1/a_81_21# -0.0191f
C103 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__a21o_1_0/X 0.00439f
C104 sky130_fd_sc_hd__a21o_1_0/a_299_297# G1 0.0137f
C105 VNB P2 0.00318f
C106 G3 sky130_fd_sc_hd__a21o_1_0/X 0.0894f
C107 VNB sky130_fd_sc_hd__a21o_1_3/a_384_47# -5.85e-20
C108 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__and4_1_0/a_303_47# 4.26e-19
C109 VNB CI 0.02f
C110 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__and4_1_0/a_27_47# 0.0588f
C111 P4 sky130_fd_sc_hd__a21o_1_2/a_299_297# 0.0108f
C112 P3 P1 0.0581f
C113 P2 sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.0301f
C114 sky130_fd_sc_hd__a21o_1_1/a_384_47# sky130_fd_sc_hd__a21o_1_1/X 4.81e-19
C115 P3 sky130_fd_sc_hd__and4_1_0/a_109_47# 0.00143f
C116 G4 P1 1.7e-20
C117 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__a21o_1_1/a_81_21# 0.00223f
C118 sky130_fd_sc_hd__a21o_1_2/X P2 0.455f
C119 G3 sky130_fd_sc_hd__a21o_1_1/a_81_21# 0.023f
C120 VPB sky130_fd_sc_hd__a21o_1_0/a_299_297# 0.00347f
C121 G3 P2 0.0287f
C122 sky130_fd_sc_hd__a21o_1_1/X sky130_fd_sc_hd__a21o_1_2/a_299_297# 0.0193f
C123 sky130_fd_sc_hd__a21o_1_2/X CI 0.00156f
C124 sky130_fd_sc_hd__and4_1_0/X sky130_fd_sc_hd__a21o_1_0/X 7.95e-21
C125 sky130_fd_sc_hd__and4_1_0/a_303_47# sky130_fd_sc_hd__and4_1_0/X 3.17e-19
C126 P4 sky130_fd_sc_hd__a21o_1_1/X 0.0428f
C127 sky130_fd_sc_hd__a21o_1_1/a_299_297# VPB -0.00193f
C128 sky130_fd_sc_hd__and4_1_0/X sky130_fd_sc_hd__and4_1_0/a_27_47# 0.00169f
C129 sky130_fd_sc_hd__and4_1_0/a_303_47# sky130_fd_sc_hd__a21o_1_0/X 5.18e-21
C130 sky130_fd_sc_hd__a21o_1_3/a_299_297# VNB -0.00378f
C131 P1 sky130_fd_sc_hd__a21o_1_3/a_81_21# 0.00196f
C132 VNB sky130_fd_sc_hd__a21o_1_0/a_384_47# -2.71e-19
C133 sky130_fd_sc_hd__and4_1_0/X P2 0.00135f
C134 VNB P1 0.0237f
C135 sky130_fd_sc_hd__and4_1_0/X sky130_fd_sc_hd__a21o_1_3/a_384_47# 7.24e-19
C136 sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__a21o_1_0/X 2.06e-20
C137 P3 sky130_fd_sc_hd__a21o_1_1/a_299_297# 0.00415f
C138 sky130_fd_sc_hd__and4_1_0/X CI 0.0308f
C139 VNB G2 0.00126f
C140 VNB sky130_fd_sc_hd__a21o_1_0/a_81_21# -0.0202f
C141 sky130_fd_sc_hd__and4_1_0/a_109_47# VNB -6.28e-20
C142 VPB sky130_fd_sc_hd__a21o_1_1/a_384_47# -4.08e-19
C143 sky130_fd_sc_hd__a21o_1_1/a_81_21# sky130_fd_sc_hd__a21o_1_0/X 0.0631f
C144 VPB sky130_fd_sc_hd__a21o_1_2/a_299_297# 0.0196f
C145 P2 sky130_fd_sc_hd__a21o_1_0/X 0.0752f
C146 sky130_fd_sc_hd__and4_1_0/a_197_47# VPB -5.24e-19
C147 P1 sky130_fd_sc_hd__a21o_1_2/a_81_21# 3.15e-20
C148 sky130_fd_sc_hd__a21o_1_1/X G1 0.00394f
C149 sky130_fd_sc_hd__a21o_1_3/a_299_297# sky130_fd_sc_hd__a21o_1_2/X 0.0173f
C150 sky130_fd_sc_hd__a21o_1_2/X P1 0.0247f
C151 P4 sky130_fd_sc_hd__a21o_1_2/a_384_47# 6.19e-21
C152 G3 P1 3.23e-21
C153 VPB P4 0.0594f
C154 sky130_fd_sc_hd__and4_1_0/a_27_47# P2 0.0709f
C155 sky130_fd_sc_hd__a21o_1_2/X G2 5.09e-20
C156 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__a21o_1_0/a_81_21# 8.44e-20
C157 P3 sky130_fd_sc_hd__a21o_1_1/a_384_47# 7.45e-20
C158 VNB sky130_fd_sc_hd__a21o_1_0/a_299_297# -0.00449f
C159 P3 sky130_fd_sc_hd__a21o_1_2/a_299_297# 0.00159f
C160 sky130_fd_sc_hd__a21o_1_2/a_384_47# sky130_fd_sc_hd__a21o_1_1/X 7.94e-20
C161 P3 sky130_fd_sc_hd__and4_1_0/a_197_47# 0.0016f
C162 sky130_fd_sc_hd__a21o_1_1/a_81_21# P2 0.0526f
C163 VPB sky130_fd_sc_hd__a21o_1_1/X 0.0255f
C164 P2 CI 2.97e-20
C165 sky130_fd_sc_hd__a21o_1_1/a_299_297# VNB -0.00449f
C166 sky130_fd_sc_hd__a21o_1_3/a_299_297# sky130_fd_sc_hd__and4_1_0/X 0.00642f
C167 P3 P4 0.2f
C168 sky130_fd_sc_hd__and4_1_0/X P1 0.00732f
C169 G4 P4 0.02f
C170 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__a21o_1_0/a_299_297# 1.65e-19
C171 sky130_fd_sc_hd__and4_1_0/a_109_47# sky130_fd_sc_hd__and4_1_0/X 1.62e-19
C172 VPB G1 0.0196f
C173 P3 sky130_fd_sc_hd__a21o_1_1/X 0.185f
C174 sky130_fd_sc_hd__a21o_1_0/a_384_47# sky130_fd_sc_hd__a21o_1_0/X 0.00135f
C175 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__a21o_1_1/a_299_297# 0.0334f
C176 P1 sky130_fd_sc_hd__a21o_1_0/X 1.23e-20
C177 G4 sky130_fd_sc_hd__a21o_1_1/X 0.0897f
C178 sky130_fd_sc_hd__a21o_1_0/X G2 0.0575f
C179 VNB sky130_fd_sc_hd__a21o_1_1/a_384_47# -1.89e-19
C180 sky130_fd_sc_hd__a21o_1_0/a_81_21# sky130_fd_sc_hd__a21o_1_0/X 0.059f
C181 sky130_fd_sc_hd__and4_1_0/a_109_47# sky130_fd_sc_hd__a21o_1_0/X 9.17e-21
C182 VPB CO -0.00363f
C183 P1 sky130_fd_sc_hd__and4_1_0/a_27_47# 0.019f
C184 VNB sky130_fd_sc_hd__a21o_1_2/a_299_297# -0.00449f
C185 sky130_fd_sc_hd__and4_1_0/a_197_47# VNB -4.52e-20
C186 VPB sky130_fd_sc_hd__a21o_1_2/a_384_47# -4.08e-19
C187 VNB P4 0.00496f
C188 sky130_fd_sc_hd__a21o_1_3/a_299_297# CI 0.00978f
C189 P1 P2 0.0215f
C190 P1 CI 2.89e-19
C191 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__a21o_1_1/a_384_47# 1.32e-20
C192 P2 G2 0.00123f
C193 sky130_fd_sc_hd__a21o_1_0/a_81_21# P2 0.00281f
C194 sky130_fd_sc_hd__and4_1_0/a_109_47# P2 2.77e-19
C195 P3 CO 0.0012f
C196 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__a21o_1_2/a_299_297# 0.0335f
C197 sky130_fd_sc_hd__a21o_1_0/X sky130_fd_sc_hd__a21o_1_0/a_299_297# 0.00259f
C198 P3 sky130_fd_sc_hd__a21o_1_2/a_384_47# 0.0013f
C199 VNB sky130_fd_sc_hd__a21o_1_1/X 0.0139f
C200 P3 VPB 0.0048f
C201 P4 sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.00149f
C202 sky130_fd_sc_hd__a21o_1_2/X P4 0.00977f
C203 G4 VPB -0.00221f
C204 VNB 0 1.71f
C205 VPB 0 4.61f
C206 sky130_fd_sc_hd__and4_1_0/X 0 0.154f
C207 P1 0 0.164f
C208 P3 0 0.297f
C209 P2 0 0.31f
C210 P4 0 0.324f
C211 sky130_fd_sc_hd__and4_1_0/a_27_47# 0 0.175f
C212 CO 0 0.0276f
C213 CI 0 0.158f
C214 sky130_fd_sc_hd__a21o_1_3/a_299_297# 0 0.0348f
C215 sky130_fd_sc_hd__a21o_1_3/a_81_21# 0 0.147f
C216 sky130_fd_sc_hd__a21o_1_2/X 0 0.168f
C217 sky130_fd_sc_hd__a21o_1_1/X 0 0.129f
C218 G4 0 0.137f
C219 sky130_fd_sc_hd__a21o_1_2/a_299_297# 0 0.0348f
C220 sky130_fd_sc_hd__a21o_1_2/a_81_21# 0 0.147f
C221 sky130_fd_sc_hd__a21o_1_0/X 0 0.223f
C222 G3 0 0.137f
C223 sky130_fd_sc_hd__a21o_1_1/a_299_297# 0 0.0348f
C224 sky130_fd_sc_hd__a21o_1_1/a_81_21# 0 0.147f
C225 G1 0 0.12f
C226 G2 0 0.163f
C227 sky130_fd_sc_hd__a21o_1_0/a_299_297# 0 0.0348f
C228 sky130_fd_sc_hd__a21o_1_0/a_81_21# 0 0.147f
.ends

.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X a_117_297# a_285_297# a_285_47#
+ a_35_297#
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.177 ps=1.69 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.138 ps=1.4 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.177 pd=1.69 as=0.177 ps=1.69 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.138 pd=1.4 as=0.0878 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.138 pd=1.4 as=0.25 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.177 pd=1.69 as=0.177 ps=1.69 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.177 pd=1.69 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.138 ps=1.4 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
C0 VGND A 0.0325f
C1 VPWR VPB 0.0689f
C2 a_117_297# B 0.00777f
C3 VGND B 0.0304f
C4 B A 0.221f
C5 VPWR X 0.0537f
C6 a_117_297# a_35_297# 0.00641f
C7 VGND a_35_297# 0.177f
C8 A a_35_297# 0.0633f
C9 VPWR a_285_47# 8.6e-19
C10 VGND VPB 0.00696f
C11 a_285_297# VPWR 0.246f
C12 A VPB 0.051f
C13 B a_35_297# 0.203f
C14 a_117_297# X 2.25e-19
C15 VGND X 0.173f
C16 B VPB 0.0697f
C17 A X 0.00166f
C18 VPB a_35_297# 0.0699f
C19 VGND a_285_47# 0.00552f
C20 B X 0.0149f
C21 VGND a_285_297# 0.00394f
C22 a_285_297# A 0.00749f
C23 X a_35_297# 0.166f
C24 B a_285_47# 3.98e-19
C25 B a_285_297# 0.0553f
C26 X VPB 0.0154f
C27 a_285_47# a_35_297# 0.00723f
C28 a_285_297# a_35_297# 0.025f
C29 a_117_297# VPWR 0.00852f
C30 VGND VPWR 0.0643f
C31 a_285_297# VPB 0.0133f
C32 VPWR A 0.0348f
C33 a_285_47# X 0.00206f
C34 a_285_297# X 0.0712f
C35 B VPWR 0.0703f
C36 VPWR a_35_297# 0.096f
C37 VGND a_117_297# 0.00177f
C38 VGND VNB 0.435f
C39 X VNB 0.0649f
C40 VPWR VNB 0.333f
C41 A VNB 0.167f
C42 B VNB 0.213f
C43 VPB VNB 0.693f
C44 a_285_297# VNB 0.00137f
C45 a_35_297# VNB 0.255f
.ends

.subckt adder_3 G1 P2 G2 G3 P4 S1 S2 S3 S4 sky130_fd_sc_hd__xor2_1_3/a_117_297# sky130_fd_sc_hd__xor2_1_3/a_35_297#
+ sky130_fd_sc_hd__a21o_1_0/a_81_21# sky130_fd_sc_hd__xor2_1_3/a_285_47# sky130_fd_sc_hd__xor2_1_0/a_285_297#
+ sky130_fd_sc_hd__a21o_1_0/a_384_47# sky130_fd_sc_hd__xor2_1_1/a_285_297# sky130_fd_sc_hd__xor2_1_0/a_35_297#
+ sky130_fd_sc_hd__xor2_1_0/a_285_47# sky130_fd_sc_hd__a21o_1_0/a_299_297# sky130_fd_sc_hd__a21o_1_1/a_81_21#
+ sky130_fd_sc_hd__xor2_1_2/a_285_297# sky130_fd_sc_hd__xor2_1_3/a_285_297# sky130_fd_sc_hd__a21o_1_1/a_299_297#
+ sky130_fd_sc_hd__a21o_1_2/a_299_297# sky130_fd_sc_hd__xor2_1_1/a_35_297# sky130_fd_sc_hd__xor2_1_3/B
+ sky130_fd_sc_hd__xor2_1_1/a_285_47# sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__a21o_1_2/a_81_21#
+ sky130_fd_sc_hd__a21o_1_2/a_384_47# sky130_fd_sc_hd__xor2_1_0/a_117_297# sky130_fd_sc_hd__xor2_1_2/a_35_297#
+ sky130_fd_sc_hd__xor2_1_2/a_285_47# sky130_fd_sc_hd__xor2_1_1/a_117_297# CI P1 SUB
+ sky130_fd_sc_hd__xor2_1_2/B sky130_fd_sc_hd__xor2_1_2/a_117_297# VPB P3
Xsky130_fd_sc_hd__xor2_1_3 P4 sky130_fd_sc_hd__xor2_1_3/B SUB SUB VPB VPB S4 sky130_fd_sc_hd__xor2_1_3/a_117_297#
+ sky130_fd_sc_hd__xor2_1_3/a_285_297# sky130_fd_sc_hd__xor2_1_3/a_285_47# sky130_fd_sc_hd__xor2_1_3/a_35_297#
+ sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__a21o_1_0 CI P1 G1 SUB SUB VPB VPB sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__a21o_1_0/a_384_47#
+ sky130_fd_sc_hd__a21o_1_0/a_81_21# sky130_fd_sc_hd__a21o_1_0/a_299_297# sky130_fd_sc_hd__a21o_1
Xsky130_fd_sc_hd__a21o_1_1 sky130_fd_sc_hd__xor2_1_1/B P2 G2 SUB SUB VPB VPB sky130_fd_sc_hd__xor2_1_2/B
+ sky130_fd_sc_hd__a21o_1_1/a_384_47# sky130_fd_sc_hd__a21o_1_1/a_81_21# sky130_fd_sc_hd__a21o_1_1/a_299_297#
+ sky130_fd_sc_hd__a21o_1
Xsky130_fd_sc_hd__a21o_1_2 sky130_fd_sc_hd__xor2_1_2/B P3 G3 SUB SUB VPB VPB sky130_fd_sc_hd__xor2_1_3/B
+ sky130_fd_sc_hd__a21o_1_2/a_384_47# sky130_fd_sc_hd__a21o_1_2/a_81_21# sky130_fd_sc_hd__a21o_1_2/a_299_297#
+ sky130_fd_sc_hd__a21o_1
Xsky130_fd_sc_hd__xor2_1_0 P1 CI SUB SUB VPB VPB S1 sky130_fd_sc_hd__xor2_1_0/a_117_297#
+ sky130_fd_sc_hd__xor2_1_0/a_285_297# sky130_fd_sc_hd__xor2_1_0/a_285_47# sky130_fd_sc_hd__xor2_1_0/a_35_297#
+ sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_1 P2 sky130_fd_sc_hd__xor2_1_1/B SUB SUB VPB VPB S2 sky130_fd_sc_hd__xor2_1_1/a_117_297#
+ sky130_fd_sc_hd__xor2_1_1/a_285_297# sky130_fd_sc_hd__xor2_1_1/a_285_47# sky130_fd_sc_hd__xor2_1_1/a_35_297#
+ sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_2 P3 sky130_fd_sc_hd__xor2_1_2/B SUB SUB VPB VPB S3 sky130_fd_sc_hd__xor2_1_2/a_117_297#
+ sky130_fd_sc_hd__xor2_1_2/a_285_297# sky130_fd_sc_hd__xor2_1_2/a_285_47# sky130_fd_sc_hd__xor2_1_2/a_35_297#
+ sky130_fd_sc_hd__xor2_1
C0 S1 S2 0.0103f
C1 sky130_fd_sc_hd__xor2_1_3/B sky130_fd_sc_hd__a21o_1_0/a_81_21# 1.96e-19
C2 P2 CI 0.186f
C3 sky130_fd_sc_hd__xor2_1_3/a_35_297# S4 0.00521f
C4 P3 sky130_fd_sc_hd__xor2_1_1/B 0.051f
C5 P3 sky130_fd_sc_hd__xor2_1_2/B 0.902f
C6 SUB sky130_fd_sc_hd__xor2_1_3/a_35_297# 0.00517f
C7 P1 sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.0139f
C8 P2 sky130_fd_sc_hd__xor2_1_1/a_285_47# 0.00118f
C9 P1 VPB 0.00988f
C10 VPB sky130_fd_sc_hd__xor2_1_1/a_285_297# 2.35e-20
C11 S3 sky130_fd_sc_hd__xor2_1_3/B 0.0617f
C12 sky130_fd_sc_hd__xor2_1_2/a_285_47# P3 0.00118f
C13 P3 S4 8.8e-19
C14 sky130_fd_sc_hd__a21o_1_0/a_81_21# sky130_fd_sc_hd__xor2_1_1/B 0.0562f
C15 P1 sky130_fd_sc_hd__a21o_1_0/a_384_47# 5.49e-19
C16 sky130_fd_sc_hd__xor2_1_0/a_285_47# P1 0.00118f
C17 sky130_fd_sc_hd__a21o_1_0/a_81_21# sky130_fd_sc_hd__xor2_1_2/B 0.00447f
C18 P1 sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.00101f
C19 P3 SUB 0.27f
C20 sky130_fd_sc_hd__xor2_1_3/B sky130_fd_sc_hd__a21o_1_1/a_384_47# 1.76e-19
C21 sky130_fd_sc_hd__xor2_1_3/a_285_47# P3 3.53e-19
C22 VPB sky130_fd_sc_hd__a21o_1_2/a_299_297# 0.0344f
C23 S1 P1 0.00593f
C24 S1 sky130_fd_sc_hd__xor2_1_1/a_285_297# 0.00137f
C25 sky130_fd_sc_hd__xor2_1_3/B sky130_fd_sc_hd__xor2_1_2/a_285_297# 0.00704f
C26 P2 sky130_fd_sc_hd__xor2_1_2/a_35_297# 6.69e-19
C27 P3 sky130_fd_sc_hd__xor2_1_3/a_35_297# 0.00203f
C28 S3 sky130_fd_sc_hd__xor2_1_1/B 3.34e-20
C29 CI G2 2.73e-19
C30 sky130_fd_sc_hd__xor2_1_0/a_117_297# VPB -2.04e-19
C31 SUB sky130_fd_sc_hd__a21o_1_0/a_81_21# -0.00347f
C32 S3 sky130_fd_sc_hd__xor2_1_2/B 0.00532f
C33 sky130_fd_sc_hd__xor2_1_3/B S2 0.0546f
C34 P1 sky130_fd_sc_hd__a21o_1_2/a_81_21# 2.85e-19
C35 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__a21o_1_0/a_299_297# 0.0526f
C36 sky130_fd_sc_hd__xor2_1_2/B sky130_fd_sc_hd__a21o_1_0/a_299_297# 0.0414f
C37 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__a21o_1_1/a_384_47# 0.00123f
C38 P2 G2 6.94e-19
C39 S1 sky130_fd_sc_hd__a21o_1_2/a_299_297# 3.56e-19
C40 sky130_fd_sc_hd__xor2_1_2/B sky130_fd_sc_hd__a21o_1_1/a_384_47# 4.32e-19
C41 S3 S4 0.0102f
C42 sky130_fd_sc_hd__a21o_1_1/a_81_21# CI 1.09e-19
C43 S3 SUB -0.00162f
C44 sky130_fd_sc_hd__xor2_1_0/a_117_297# S1 4.28e-19
C45 S2 sky130_fd_sc_hd__xor2_1_1/B 0.00554f
C46 SUB sky130_fd_sc_hd__a21o_1_0/a_299_297# -0.00435f
C47 sky130_fd_sc_hd__xor2_1_2/B S2 0.00962f
C48 sky130_fd_sc_hd__a21o_1_1/a_81_21# P2 0.00611f
C49 S3 sky130_fd_sc_hd__xor2_1_3/a_35_297# 0.0518f
C50 SUB sky130_fd_sc_hd__xor2_1_2/a_285_297# -0.00394f
C51 P1 sky130_fd_sc_hd__xor2_1_3/B 0.0733f
C52 sky130_fd_sc_hd__xor2_1_3/B sky130_fd_sc_hd__xor2_1_1/a_285_297# 0.00704f
C53 SUB S2 -0.00162f
C54 sky130_fd_sc_hd__xor2_1_0/a_35_297# CI 0.0235f
C55 CI VPB 0.00219f
C56 P3 S3 0.00706f
C57 VPB sky130_fd_sc_hd__xor2_1_1/a_117_297# 2.29e-20
C58 CI sky130_fd_sc_hd__a21o_1_0/a_384_47# 0.00162f
C59 sky130_fd_sc_hd__xor2_1_0/a_35_297# P2 0.00129f
C60 sky130_fd_sc_hd__a21o_1_2/a_299_297# sky130_fd_sc_hd__xor2_1_3/B 6.06e-19
C61 CI sky130_fd_sc_hd__xor2_1_1/a_35_297# 7.26e-21
C62 P4 VPB 0.0224f
C63 P2 VPB 0.0257f
C64 P1 sky130_fd_sc_hd__xor2_1_1/B 0.132f
C65 P2 sky130_fd_sc_hd__a21o_1_1/a_299_297# 0.00664f
C66 VPB sky130_fd_sc_hd__xor2_1_1/a_285_47# -7.24e-19
C67 P1 sky130_fd_sc_hd__xor2_1_2/B 0.183f
C68 sky130_fd_sc_hd__xor2_1_2/a_117_297# VPB 2.25e-20
C69 S1 CI 0.002f
C70 sky130_fd_sc_hd__xor2_1_0/a_285_47# P2 4.62e-19
C71 sky130_fd_sc_hd__a21o_1_1/a_81_21# G2 0.0275f
C72 P2 sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.0178f
C73 P1 G3 6.62e-19
C74 S1 sky130_fd_sc_hd__xor2_1_1/a_117_297# 0.00102f
C75 P3 S2 0.00112f
C76 CI sky130_fd_sc_hd__a21o_1_2/a_81_21# 1.2e-19
C77 sky130_fd_sc_hd__a21o_1_2/a_299_297# sky130_fd_sc_hd__xor2_1_1/B 0.0519f
C78 S1 P2 0.00354f
C79 sky130_fd_sc_hd__a21o_1_2/a_299_297# sky130_fd_sc_hd__xor2_1_2/B 0.00554f
C80 P1 SUB 1f
C81 CI G1 0.0805f
C82 SUB sky130_fd_sc_hd__xor2_1_1/a_285_297# -0.00394f
C83 S1 sky130_fd_sc_hd__xor2_1_2/a_117_297# 2.46e-20
C84 sky130_fd_sc_hd__xor2_1_0/a_117_297# sky130_fd_sc_hd__xor2_1_1/B 0.00427f
C85 VPB sky130_fd_sc_hd__xor2_1_2/a_35_297# 0.00796f
C86 P2 sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.0197f
C87 sky130_fd_sc_hd__xor2_1_0/a_117_297# sky130_fd_sc_hd__xor2_1_2/B 2.27e-19
C88 sky130_fd_sc_hd__xor2_1_2/a_35_297# sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.00123f
C89 sky130_fd_sc_hd__a21o_1_2/a_299_297# SUB -0.00449f
C90 VPB G2 0.00129f
C91 S3 sky130_fd_sc_hd__xor2_1_2/a_285_297# 0.00453f
C92 S1 sky130_fd_sc_hd__xor2_1_2/a_35_297# 2.99e-20
C93 sky130_fd_sc_hd__xor2_1_0/a_117_297# SUB -0.00177f
C94 sky130_fd_sc_hd__xor2_1_3/a_285_297# S4 0.00453f
C95 S3 S2 0.0102f
C96 P1 P3 0.0282f
C97 CI sky130_fd_sc_hd__xor2_1_3/B 0.0784f
C98 sky130_fd_sc_hd__a21o_1_1/a_81_21# VPB -0.00424f
C99 sky130_fd_sc_hd__xor2_1_1/a_117_297# sky130_fd_sc_hd__xor2_1_3/B 0.00134f
C100 P4 sky130_fd_sc_hd__xor2_1_3/B 0.104f
C101 P2 sky130_fd_sc_hd__xor2_1_3/B 0.107f
C102 sky130_fd_sc_hd__xor2_1_0/a_35_297# sky130_fd_sc_hd__a21o_1_2/a_384_47# 6.06e-21
C103 S2 sky130_fd_sc_hd__xor2_1_2/a_285_297# 0.00111f
C104 sky130_fd_sc_hd__xor2_1_3/B sky130_fd_sc_hd__xor2_1_1/a_285_47# 0.00253f
C105 P1 sky130_fd_sc_hd__a21o_1_0/a_81_21# 7.84e-20
C106 P3 sky130_fd_sc_hd__a21o_1_2/a_299_297# 0.00623f
C107 VPB sky130_fd_sc_hd__a21o_1_2/a_384_47# -4.08e-19
C108 sky130_fd_sc_hd__xor2_1_2/a_117_297# sky130_fd_sc_hd__xor2_1_3/B 0.00134f
C109 CI sky130_fd_sc_hd__xor2_1_1/B 0.155f
C110 G2 G1 1.42e-20
C111 CI sky130_fd_sc_hd__xor2_1_2/B 0.818f
C112 sky130_fd_sc_hd__xor2_1_1/a_117_297# sky130_fd_sc_hd__xor2_1_1/B 0.00269f
C113 CI G3 2.35e-19
C114 sky130_fd_sc_hd__xor2_1_0/a_35_297# VPB 0.042f
C115 P4 sky130_fd_sc_hd__xor2_1_1/B 9.9e-21
C116 P2 sky130_fd_sc_hd__xor2_1_1/B 0.223f
C117 S3 sky130_fd_sc_hd__xor2_1_1/a_285_297# 8.64e-20
C118 P2 sky130_fd_sc_hd__xor2_1_2/B 0.163f
C119 VPB sky130_fd_sc_hd__a21o_1_1/a_299_297# 0.0016f
C120 VPB sky130_fd_sc_hd__xor2_1_0/a_285_297# -3.91e-19
C121 sky130_fd_sc_hd__xor2_1_1/a_285_47# sky130_fd_sc_hd__xor2_1_2/B 5.8e-19
C122 sky130_fd_sc_hd__xor2_1_2/a_35_297# sky130_fd_sc_hd__xor2_1_3/B 0.0908f
C123 P1 sky130_fd_sc_hd__a21o_1_0/a_299_297# 0.00669f
C124 sky130_fd_sc_hd__xor2_1_2/a_117_297# sky130_fd_sc_hd__xor2_1_2/B 0.00267f
C125 CI SUB 0.176f
C126 sky130_fd_sc_hd__xor2_1_0/a_35_297# sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.00128f
C127 VPB sky130_fd_sc_hd__a21o_1_0/a_384_47# -4.08e-19
C128 sky130_fd_sc_hd__xor2_1_0/a_285_47# VPB -8.6e-19
C129 P2 G3 0.0223f
C130 VPB sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.00693f
C131 sky130_fd_sc_hd__xor2_1_1/a_117_297# SUB -0.00177f
C132 P4 S4 0.00239f
C133 S1 sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.00396f
C134 sky130_fd_sc_hd__xor2_1_3/B G2 2.64e-19
C135 P4 SUB 0.0233f
C136 P2 SUB 0.384f
C137 sky130_fd_sc_hd__xor2_1_3/a_117_297# VPB 2.25e-20
C138 S1 VPB 0.0368f
C139 SUB sky130_fd_sc_hd__xor2_1_1/a_285_47# -4.65e-19
C140 S1 sky130_fd_sc_hd__a21o_1_1/a_299_297# 8.32e-20
C141 S1 sky130_fd_sc_hd__xor2_1_0/a_285_297# 0.00385f
C142 sky130_fd_sc_hd__xor2_1_2/a_117_297# SUB -0.00177f
C143 S2 sky130_fd_sc_hd__xor2_1_1/a_285_297# 0.00293f
C144 sky130_fd_sc_hd__xor2_1_0/a_35_297# sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.00109f
C145 sky130_fd_sc_hd__xor2_1_2/a_35_297# sky130_fd_sc_hd__xor2_1_1/B 6.93e-20
C146 VPB sky130_fd_sc_hd__a21o_1_2/a_81_21# -0.00306f
C147 sky130_fd_sc_hd__xor2_1_2/a_35_297# sky130_fd_sc_hd__xor2_1_2/B 0.0262f
C148 S3 sky130_fd_sc_hd__xor2_1_3/a_285_297# 0.00135f
C149 S1 sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.0535f
C150 P4 sky130_fd_sc_hd__xor2_1_3/a_35_297# 0.0132f
C151 P2 sky130_fd_sc_hd__xor2_1_3/a_35_297# 3.67e-21
C152 sky130_fd_sc_hd__a21o_1_1/a_81_21# sky130_fd_sc_hd__xor2_1_3/B 0.00303f
C153 VPB G1 0.00163f
C154 P3 CI 0.346f
C155 G2 sky130_fd_sc_hd__xor2_1_1/B 0.13f
C156 sky130_fd_sc_hd__xor2_1_2/B G2 0.0266f
C157 sky130_fd_sc_hd__xor2_1_2/a_35_297# SUB -0.0113f
C158 sky130_fd_sc_hd__xor2_1_3/B sky130_fd_sc_hd__a21o_1_2/a_384_47# 0.00131f
C159 S1 sky130_fd_sc_hd__a21o_1_2/a_81_21# 2.24e-19
C160 P4 P3 4.73e-19
C161 P3 P2 0.608f
C162 CI sky130_fd_sc_hd__a21o_1_0/a_81_21# 0.0177f
C163 sky130_fd_sc_hd__a21o_1_1/a_81_21# sky130_fd_sc_hd__xor2_1_1/B 0.0601f
C164 sky130_fd_sc_hd__a21o_1_1/a_81_21# sky130_fd_sc_hd__xor2_1_2/B 0.0211f
C165 SUB G2 0.0237f
C166 sky130_fd_sc_hd__xor2_1_2/a_35_297# sky130_fd_sc_hd__xor2_1_3/a_35_297# 0.00123f
C167 sky130_fd_sc_hd__xor2_1_0/a_35_297# sky130_fd_sc_hd__xor2_1_3/B 0.0707f
C168 VPB sky130_fd_sc_hd__xor2_1_3/B 0.167f
C169 sky130_fd_sc_hd__xor2_1_3/B sky130_fd_sc_hd__a21o_1_1/a_299_297# 0.0322f
C170 sky130_fd_sc_hd__xor2_1_3/B sky130_fd_sc_hd__xor2_1_0/a_285_297# 1.77e-19
C171 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__a21o_1_2/a_384_47# 2.81e-20
C172 sky130_fd_sc_hd__xor2_1_2/B sky130_fd_sc_hd__a21o_1_2/a_384_47# 0.00105f
C173 sky130_fd_sc_hd__xor2_1_3/B sky130_fd_sc_hd__a21o_1_0/a_384_47# 2.82e-20
C174 sky130_fd_sc_hd__xor2_1_0/a_285_47# sky130_fd_sc_hd__xor2_1_3/B 0.00255f
C175 sky130_fd_sc_hd__xor2_1_1/a_117_297# S3 1.88e-20
C176 sky130_fd_sc_hd__xor2_1_3/B sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.0714f
C177 sky130_fd_sc_hd__a21o_1_1/a_81_21# SUB -0.00243f
C178 P3 sky130_fd_sc_hd__xor2_1_2/a_35_297# 0.0152f
C179 CI sky130_fd_sc_hd__a21o_1_0/a_299_297# 0.00517f
C180 P4 S3 0.00111f
C181 sky130_fd_sc_hd__xor2_1_0/a_35_297# sky130_fd_sc_hd__xor2_1_1/B 0.0678f
C182 P2 S3 2.48e-20
C183 sky130_fd_sc_hd__xor2_1_3/a_117_297# sky130_fd_sc_hd__xor2_1_3/B 0.00267f
C184 S1 sky130_fd_sc_hd__xor2_1_3/B 0.0317f
C185 sky130_fd_sc_hd__xor2_1_0/a_35_297# sky130_fd_sc_hd__xor2_1_2/B 0.00271f
C186 VPB sky130_fd_sc_hd__xor2_1_1/B 0.743f
C187 SUB sky130_fd_sc_hd__a21o_1_2/a_384_47# -2.27e-19
C188 sky130_fd_sc_hd__xor2_1_2/a_117_297# S3 6.67e-19
C189 sky130_fd_sc_hd__a21o_1_1/a_299_297# sky130_fd_sc_hd__xor2_1_1/B 0.0587f
C190 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__xor2_1_0/a_285_297# 0.036f
C191 VPB sky130_fd_sc_hd__xor2_1_2/B 0.108f
C192 sky130_fd_sc_hd__xor2_1_2/B sky130_fd_sc_hd__a21o_1_1/a_299_297# 0.00516f
C193 sky130_fd_sc_hd__xor2_1_3/B sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.0563f
C194 sky130_fd_sc_hd__xor2_1_0/a_35_297# G3 6.72e-20
C195 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__a21o_1_0/a_384_47# 3.85e-19
C196 P2 sky130_fd_sc_hd__a21o_1_1/a_384_47# 6.47e-19
C197 sky130_fd_sc_hd__xor2_1_0/a_285_47# sky130_fd_sc_hd__xor2_1_1/B 2.47e-19
C198 sky130_fd_sc_hd__xor2_1_2/B sky130_fd_sc_hd__a21o_1_0/a_384_47# 1.35e-20
C199 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.0394f
C200 VPB G3 0.00152f
C201 sky130_fd_sc_hd__xor2_1_3/B G1 1.88e-20
C202 sky130_fd_sc_hd__xor2_1_1/a_117_297# S2 5.82e-19
C203 sky130_fd_sc_hd__xor2_1_2/B sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.0151f
C204 sky130_fd_sc_hd__xor2_1_2/a_285_47# VPB -7.24e-19
C205 VPB S4 0.0296f
C206 sky130_fd_sc_hd__xor2_1_0/a_35_297# SUB -0.0143f
C207 sky130_fd_sc_hd__a21o_1_0/a_81_21# G2 1.77e-20
C208 S1 sky130_fd_sc_hd__xor2_1_1/B 0.112f
C209 P2 S2 0.0068f
C210 VPB SUB -0.376f
C211 S1 sky130_fd_sc_hd__xor2_1_2/B 1.38e-19
C212 SUB sky130_fd_sc_hd__a21o_1_1/a_299_297# -0.00436f
C213 SUB sky130_fd_sc_hd__xor2_1_0/a_285_297# -0.00394f
C214 sky130_fd_sc_hd__xor2_1_2/a_35_297# S3 0.00495f
C215 sky130_fd_sc_hd__xor2_1_2/a_117_297# S2 8.82e-19
C216 sky130_fd_sc_hd__a21o_1_2/a_81_21# sky130_fd_sc_hd__xor2_1_1/B 0.0491f
C217 SUB sky130_fd_sc_hd__a21o_1_0/a_384_47# 4.44e-34
C218 sky130_fd_sc_hd__xor2_1_0/a_285_47# SUB -4.65e-19
C219 sky130_fd_sc_hd__xor2_1_2/B sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.0116f
C220 S1 G3 8.29e-20
C221 SUB sky130_fd_sc_hd__xor2_1_1/a_35_297# -0.0109f
C222 P3 sky130_fd_sc_hd__a21o_1_2/a_384_47# 5.7e-19
C223 VPB sky130_fd_sc_hd__xor2_1_3/a_35_297# 0.00512f
C224 sky130_fd_sc_hd__xor2_1_1/B G1 0.0614f
C225 sky130_fd_sc_hd__xor2_1_3/a_117_297# S4 6.67e-19
C226 sky130_fd_sc_hd__xor2_1_2/B G1 0.0014f
C227 G3 sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.0232f
C228 sky130_fd_sc_hd__xor2_1_3/a_117_297# SUB -8.18e-19
C229 S1 SUB -0.00328f
C230 P1 CI 0.544f
C231 sky130_fd_sc_hd__xor2_1_0/a_35_297# P3 0.00793f
C232 SUB sky130_fd_sc_hd__a21o_1_2/a_81_21# -0.0181f
C233 sky130_fd_sc_hd__xor2_1_2/a_35_297# S2 0.0515f
C234 P3 VPB 0.0315f
C235 SUB G1 0.023f
C236 P1 P2 0.6f
C237 P3 sky130_fd_sc_hd__xor2_1_1/a_35_297# 2.02e-19
C238 sky130_fd_sc_hd__xor2_1_3/B sky130_fd_sc_hd__xor2_1_1/B 0.398f
C239 VPB sky130_fd_sc_hd__a21o_1_0/a_81_21# -0.00793f
C240 sky130_fd_sc_hd__xor2_1_3/B sky130_fd_sc_hd__xor2_1_2/B 0.171f
C241 S1 P3 2.04e-19
C242 sky130_fd_sc_hd__xor2_1_0/a_117_297# CI 9.44e-19
C243 G3 sky130_fd_sc_hd__xor2_1_3/B 0.0517f
C244 P3 sky130_fd_sc_hd__a21o_1_2/a_81_21# 4.57e-20
C245 sky130_fd_sc_hd__xor2_1_2/a_285_47# sky130_fd_sc_hd__xor2_1_3/B 0.00259f
C246 sky130_fd_sc_hd__xor2_1_3/B S4 0.00601f
C247 VPB S3 0.041f
C248 SUB sky130_fd_sc_hd__xor2_1_3/B 1.3f
C249 sky130_fd_sc_hd__xor2_1_2/B sky130_fd_sc_hd__xor2_1_1/B 0.161f
C250 sky130_fd_sc_hd__xor2_1_3/a_285_47# sky130_fd_sc_hd__xor2_1_3/B 3.65e-19
C251 VPB sky130_fd_sc_hd__a21o_1_0/a_299_297# 0.0016f
C252 S3 sky130_fd_sc_hd__xor2_1_1/a_35_297# 3.35e-20
C253 VPB sky130_fd_sc_hd__a21o_1_1/a_384_47# -4.08e-19
C254 G3 sky130_fd_sc_hd__xor2_1_1/B 0.0538f
C255 P1 G2 0.0104f
C256 sky130_fd_sc_hd__xor2_1_3/B sky130_fd_sc_hd__xor2_1_3/a_35_297# 0.0593f
C257 G3 sky130_fd_sc_hd__xor2_1_2/B 0.0811f
C258 sky130_fd_sc_hd__a21o_1_0/a_81_21# G1 0.0272f
C259 VPB sky130_fd_sc_hd__xor2_1_2/a_285_297# 2.35e-20
C260 sky130_fd_sc_hd__xor2_1_3/a_117_297# S3 0.00101f
C261 S1 S3 3.29e-19
C262 SUB sky130_fd_sc_hd__xor2_1_1/B 0.137f
C263 VPB S2 0.0397f
C264 SUB sky130_fd_sc_hd__xor2_1_2/B 0.233f
C265 P3 sky130_fd_sc_hd__xor2_1_3/B 0.159f
C266 sky130_fd_sc_hd__a21o_1_1/a_81_21# P1 0.0152f
C267 SUB G3 8.34e-19
C268 sky130_fd_sc_hd__xor2_1_3/a_35_297# sky130_fd_sc_hd__xor2_1_1/B 5.05e-21
C269 S2 sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.00476f
C270 sky130_fd_sc_hd__xor2_1_2/a_285_47# SUB -4.65e-19
C271 S1 sky130_fd_sc_hd__xor2_1_2/a_285_297# 4.46e-20
C272 SUB S4 0.0195f
C273 S3 0 0.0366f
C274 P3 0 0.733f
C275 sky130_fd_sc_hd__xor2_1_2/a_285_297# 0 0.00137f
C276 sky130_fd_sc_hd__xor2_1_2/a_35_297# 0 0.255f
C277 SUB 0 1.99f
C278 S2 0 0.0353f
C279 P2 0 0.625f
C280 sky130_fd_sc_hd__xor2_1_1/B 0 0.486f
C281 VPB 0 6.64f
C282 sky130_fd_sc_hd__xor2_1_1/a_285_297# 0 0.00137f
C283 sky130_fd_sc_hd__xor2_1_1/a_35_297# 0 0.255f
C284 S1 0 0.0372f
C285 P1 0 0.561f
C286 CI 0 0.811f
C287 sky130_fd_sc_hd__xor2_1_0/a_285_297# 0 0.00137f
C288 sky130_fd_sc_hd__xor2_1_0/a_35_297# 0 0.255f
C289 sky130_fd_sc_hd__xor2_1_3/B 0 0.336f
C290 sky130_fd_sc_hd__xor2_1_2/B 0 1.53f
C291 G3 0 0.135f
C292 sky130_fd_sc_hd__a21o_1_2/a_299_297# 0 0.0348f
C293 sky130_fd_sc_hd__a21o_1_2/a_81_21# 0 0.147f
C294 G2 0 0.134f
C295 sky130_fd_sc_hd__a21o_1_1/a_299_297# 0 0.0348f
C296 sky130_fd_sc_hd__a21o_1_1/a_81_21# 0 0.147f
C297 G1 0 0.156f
C298 sky130_fd_sc_hd__a21o_1_0/a_299_297# 0 0.0348f
C299 sky130_fd_sc_hd__a21o_1_0/a_81_21# 0 0.147f
C300 S4 0 0.113f
C301 P4 0 0.21f
C302 sky130_fd_sc_hd__xor2_1_3/a_285_297# 0 0.00137f
C303 sky130_fd_sc_hd__xor2_1_3/a_35_297# 0 0.255f
.ends

.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X a_145_75# a_59_75#
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.103 pd=0.954 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.245 ps=2.27 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.816 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.103 ps=0.954 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.136 ps=1.26 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
C0 VPB X 0.0127f
C1 a_145_75# VPWR 6.31e-19
C2 VGND A 0.0147f
C3 B X 0.00276f
C4 a_59_75# A 0.0809f
C5 VPB B 0.0629f
C6 a_59_75# VGND 0.116f
C7 VPWR A 0.0362f
C8 VPWR VGND 0.0461f
C9 VPWR a_59_75# 0.15f
C10 a_145_75# X 5.76e-19
C11 A X 1.68e-19
C12 VGND X 0.0993f
C13 VPB A 0.0806f
C14 a_59_75# X 0.109f
C15 VPB VGND 0.008f
C16 VPB a_59_75# 0.0563f
C17 A B 0.0971f
C18 VPWR X 0.111f
C19 VGND B 0.0115f
C20 VPB VPWR 0.0729f
C21 a_59_75# B 0.143f
C22 VPWR B 0.0117f
C23 a_145_75# VGND 0.00468f
C24 a_145_75# a_59_75# 0.00658f
C25 VGND VNB 0.311f
C26 X VNB 0.1f
C27 B VNB 0.113f
C28 A VNB 0.174f
C29 VPWR VNB 0.273f
C30 VPB VNB 0.516f
C31 a_59_75# VNB 0.177f
.ends

.subckt adder_1 A1 B1 A2 B2 A3 B3 A4 B4 G1 P1 G2 P2 G3 P3 G4 P4 sky130_fd_sc_hd__xor2_1_3/a_117_297#
+ sky130_fd_sc_hd__xor2_1_3/a_35_297# sky130_fd_sc_hd__xor2_1_3/a_285_47# sky130_fd_sc_hd__and2_1_3/a_145_75#
+ sky130_fd_sc_hd__and2_1_2/a_59_75# sky130_fd_sc_hd__xor2_1_0/a_285_297# sky130_fd_sc_hd__xor2_1_1/a_285_297#
+ sky130_fd_sc_hd__xor2_1_0/a_35_297# sky130_fd_sc_hd__xor2_1_0/a_285_47# sky130_fd_sc_hd__xor2_1_2/a_285_297#
+ sky130_fd_sc_hd__and2_1_0/a_145_75# sky130_fd_sc_hd__xor2_1_3/a_285_297# sky130_fd_sc_hd__and2_1_3/a_59_75#
+ sky130_fd_sc_hd__xor2_1_1/a_35_297# sky130_fd_sc_hd__xor2_1_1/a_285_47# sky130_fd_sc_hd__and2_1_1/a_145_75#
+ sky130_fd_sc_hd__and2_1_0/a_59_75# sky130_fd_sc_hd__xor2_1_0/a_117_297# sky130_fd_sc_hd__xor2_1_2/a_35_297#
+ sky130_fd_sc_hd__xor2_1_2/a_285_47# sky130_fd_sc_hd__xor2_1_1/a_117_297# sky130_fd_sc_hd__and2_1_2/a_145_75#
+ SUB sky130_fd_sc_hd__and2_1_1/a_59_75# sky130_fd_sc_hd__xor2_1_2/a_117_297# VDD
Xsky130_fd_sc_hd__xor2_1_3 A4 B4 SUB SUB VDD VDD P4 sky130_fd_sc_hd__xor2_1_3/a_117_297#
+ sky130_fd_sc_hd__xor2_1_3/a_285_297# sky130_fd_sc_hd__xor2_1_3/a_285_47# sky130_fd_sc_hd__xor2_1_3/a_35_297#
+ sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__and2_1_0 A1 B1 SUB SUB VDD VDD G1 sky130_fd_sc_hd__and2_1_0/a_145_75#
+ sky130_fd_sc_hd__and2_1_0/a_59_75# sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__and2_1_1 A2 B2 SUB SUB VDD VDD G2 sky130_fd_sc_hd__and2_1_1/a_145_75#
+ sky130_fd_sc_hd__and2_1_1/a_59_75# sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__and2_1_2 A3 B3 SUB SUB VDD VDD G3 sky130_fd_sc_hd__and2_1_2/a_145_75#
+ sky130_fd_sc_hd__and2_1_2/a_59_75# sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__and2_1_3 A4 B4 SUB SUB VDD VDD G4 sky130_fd_sc_hd__and2_1_3/a_145_75#
+ sky130_fd_sc_hd__and2_1_3/a_59_75# sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__xor2_1_0 A1 B1 SUB SUB VDD VDD P1 sky130_fd_sc_hd__xor2_1_0/a_117_297#
+ sky130_fd_sc_hd__xor2_1_0/a_285_297# sky130_fd_sc_hd__xor2_1_0/a_285_47# sky130_fd_sc_hd__xor2_1_0/a_35_297#
+ sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_1 A2 B2 SUB SUB VDD VDD P2 sky130_fd_sc_hd__xor2_1_1/a_117_297#
+ sky130_fd_sc_hd__xor2_1_1/a_285_297# sky130_fd_sc_hd__xor2_1_1/a_285_47# sky130_fd_sc_hd__xor2_1_1/a_35_297#
+ sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_2 A3 B3 SUB SUB VDD VDD P3 sky130_fd_sc_hd__xor2_1_2/a_117_297#
+ sky130_fd_sc_hd__xor2_1_2/a_285_297# sky130_fd_sc_hd__xor2_1_2/a_285_47# sky130_fd_sc_hd__xor2_1_2/a_35_297#
+ sky130_fd_sc_hd__xor2_1
C0 B3 sky130_fd_sc_hd__and2_1_3/a_59_75# 4.1e-19
C1 sky130_fd_sc_hd__xor2_1_2/a_117_297# P3 2.16e-19
C2 sky130_fd_sc_hd__xor2_1_3/a_117_297# G4 7.98e-19
C3 B2 sky130_fd_sc_hd__and2_1_0/a_145_75# 1.12e-21
C4 A2 SUB 0.0431f
C5 P2 SUB 0.00985f
C6 B4 sky130_fd_sc_hd__and2_1_3/a_59_75# 0.0576f
C7 A2 sky130_fd_sc_hd__and2_1_1/a_145_75# 0.00119f
C8 A1 G1 0.0701f
C9 sky130_fd_sc_hd__xor2_1_3/a_35_297# B4 0.0414f
C10 sky130_fd_sc_hd__xor2_1_3/a_285_297# A4 6.41e-19
C11 G3 A4 1.39e-19
C12 sky130_fd_sc_hd__xor2_1_0/a_285_297# G1 5.75e-19
C13 sky130_fd_sc_hd__xor2_1_2/a_35_297# sky130_fd_sc_hd__and2_1_3/a_59_75# 0.00179f
C14 B3 B4 0.00433f
C15 sky130_fd_sc_hd__and2_1_2/a_145_75# A3 0.00119f
C16 B3 sky130_fd_sc_hd__xor2_1_2/a_35_297# 0.0715f
C17 sky130_fd_sc_hd__xor2_1_2/a_117_297# A3 0.00414f
C18 A1 SUB 0.0438f
C19 A2 VDD 0.198f
C20 VDD P2 0.0747f
C21 A2 B1 0.00281f
C22 sky130_fd_sc_hd__xor2_1_2/a_285_47# SUB -2.55e-19
C23 B2 P1 8.23e-19
C24 A2 G2 0.071f
C25 P2 G2 0.00318f
C26 B4 sky130_fd_sc_hd__xor2_1_2/a_35_297# 4.2e-19
C27 sky130_fd_sc_hd__xor2_1_2/a_117_297# G4 1.25e-19
C28 sky130_fd_sc_hd__xor2_1_3/a_117_297# A4 0.00414f
C29 P1 sky130_fd_sc_hd__and2_1_0/a_59_75# 1.33e-19
C30 B2 sky130_fd_sc_hd__and2_1_2/a_59_75# 1.27e-19
C31 B2 sky130_fd_sc_hd__xor2_1_1/a_285_297# 1.19e-19
C32 sky130_fd_sc_hd__and2_1_1/a_59_75# P1 0.00746f
C33 G3 sky130_fd_sc_hd__xor2_1_3/a_117_297# 9e-22
C34 B2 G1 7.99e-20
C35 VDD A1 0.182f
C36 A1 B1 0.264f
C37 VDD sky130_fd_sc_hd__xor2_1_2/a_285_47# -8.2e-19
C38 sky130_fd_sc_hd__xor2_1_0/a_285_297# VDD 4.65e-20
C39 G1 sky130_fd_sc_hd__and2_1_0/a_59_75# 0.00228f
C40 A1 G2 1.14e-19
C41 B3 A2 1e-19
C42 sky130_fd_sc_hd__xor2_1_0/a_285_297# B1 1.19e-19
C43 B3 P2 5.55e-19
C44 P3 sky130_fd_sc_hd__and2_1_2/a_59_75# 9.47e-20
C45 sky130_fd_sc_hd__xor2_1_0/a_285_297# G2 3.25e-19
C46 B2 SUB 0.157f
C47 sky130_fd_sc_hd__and2_1_1/a_59_75# G1 8.11e-20
C48 P3 sky130_fd_sc_hd__xor2_1_1/a_285_297# 2.3e-20
C49 B2 sky130_fd_sc_hd__and2_1_1/a_145_75# 2.28e-20
C50 sky130_fd_sc_hd__and2_1_0/a_59_75# SUB -0.00661f
C51 P2 sky130_fd_sc_hd__xor2_1_2/a_35_297# 1.96e-20
C52 P1 A3 1.12e-21
C53 sky130_fd_sc_hd__and2_1_1/a_59_75# SUB 0.00649f
C54 B3 sky130_fd_sc_hd__xor2_1_2/a_285_47# 0.00257f
C55 P4 SUB 0.00985f
C56 P3 SUB 0.0125f
C57 A3 sky130_fd_sc_hd__and2_1_2/a_59_75# 0.0594f
C58 G3 sky130_fd_sc_hd__xor2_1_2/a_117_297# 7.99e-19
C59 B2 VDD 0.00698f
C60 B2 B1 0.00218f
C61 VDD sky130_fd_sc_hd__and2_1_0/a_59_75# -0.00241f
C62 A3 sky130_fd_sc_hd__xor2_1_1/a_285_297# 4.35e-19
C63 B2 G2 0.042f
C64 B1 sky130_fd_sc_hd__and2_1_0/a_59_75# 0.0544f
C65 B3 sky130_fd_sc_hd__xor2_1_1/a_285_47# 3.82e-20
C66 B4 sky130_fd_sc_hd__xor2_1_3/a_285_47# 2.19e-19
C67 sky130_fd_sc_hd__and2_1_1/a_59_75# VDD -7.45e-19
C68 sky130_fd_sc_hd__and2_1_1/a_59_75# B1 9.42e-20
C69 VDD P4 0.0238f
C70 A2 P2 0.00233f
C71 VDD P3 0.0448f
C72 sky130_fd_sc_hd__and2_1_1/a_59_75# G2 0.00228f
C73 sky130_fd_sc_hd__xor2_1_2/a_285_297# SUB -0.00166f
C74 A3 SUB 0.0164f
C75 B3 B2 0.00271f
C76 G4 SUB -1.95e-19
C77 P4 sky130_fd_sc_hd__and2_1_3/a_59_75# 2.68e-20
C78 A2 A1 0.00698f
C79 P3 sky130_fd_sc_hd__and2_1_3/a_59_75# 0.00722f
C80 A1 P2 1.59e-21
C81 sky130_fd_sc_hd__xor2_1_3/a_35_297# P4 0.00234f
C82 sky130_fd_sc_hd__xor2_1_0/a_285_297# A2 3.31e-19
C83 sky130_fd_sc_hd__xor2_1_0/a_285_297# P2 1.01e-20
C84 sky130_fd_sc_hd__xor2_1_3/a_35_297# P3 1.05e-19
C85 sky130_fd_sc_hd__xor2_1_0/a_285_47# B1 2.19e-19
C86 VDD sky130_fd_sc_hd__xor2_1_2/a_285_297# 4.65e-20
C87 A4 sky130_fd_sc_hd__and2_1_2/a_59_75# 4.2e-20
C88 VDD A3 0.208f
C89 B3 P3 0.00724f
C90 G2 A3 6.19e-20
C91 B4 P4 0.00126f
C92 P3 B4 7.42e-19
C93 VDD G4 0.0395f
C94 G3 sky130_fd_sc_hd__and2_1_2/a_59_75# 0.0029f
C95 sky130_fd_sc_hd__xor2_1_0/a_35_297# P1 0.00153f
C96 sky130_fd_sc_hd__xor2_1_2/a_35_297# P4 5.81e-21
C97 sky130_fd_sc_hd__xor2_1_0/a_285_297# A1 6.41e-19
C98 P3 sky130_fd_sc_hd__xor2_1_2/a_35_297# 0.00192f
C99 sky130_fd_sc_hd__xor2_1_1/a_35_297# P1 1.51e-19
C100 A4 SUB 0.0446f
C101 B3 sky130_fd_sc_hd__xor2_1_2/a_285_297# 0.00523f
C102 B3 A3 0.294f
C103 sky130_fd_sc_hd__xor2_1_0/a_117_297# P1 3.4e-19
C104 sky130_fd_sc_hd__xor2_1_1/a_35_297# sky130_fd_sc_hd__and2_1_2/a_59_75# 0.00133f
C105 A2 B2 0.256f
C106 G4 sky130_fd_sc_hd__and2_1_3/a_59_75# 0.0026f
C107 B2 P2 0.00129f
C108 sky130_fd_sc_hd__xor2_1_0/a_35_297# G1 0.0663f
C109 sky130_fd_sc_hd__xor2_1_3/a_35_297# G4 0.0665f
C110 A2 sky130_fd_sc_hd__and2_1_0/a_59_75# 4.2e-20
C111 G3 SUB -1.95e-19
C112 B3 G4 9.35e-20
C113 A2 sky130_fd_sc_hd__and2_1_1/a_59_75# 0.0589f
C114 A3 sky130_fd_sc_hd__xor2_1_2/a_35_297# 0.0336f
C115 A4 sky130_fd_sc_hd__and2_1_3/a_145_75# 0.00119f
C116 sky130_fd_sc_hd__xor2_1_0/a_35_297# SUB -0.00339f
C117 sky130_fd_sc_hd__xor2_1_0/a_117_297# G1 7.26e-19
C118 sky130_fd_sc_hd__and2_1_1/a_59_75# P2 4.05e-20
C119 VDD A4 0.197f
C120 B4 G4 0.0423f
C121 P2 P3 2.24e-20
C122 B2 A1 1.47e-19
C123 sky130_fd_sc_hd__xor2_1_1/a_35_297# SUB -0.00565f
C124 G4 sky130_fd_sc_hd__xor2_1_2/a_35_297# 2.26e-19
C125 A1 sky130_fd_sc_hd__and2_1_0/a_59_75# 0.0581f
C126 sky130_fd_sc_hd__xor2_1_3/a_117_297# SUB -0.00177f
C127 sky130_fd_sc_hd__xor2_1_3/a_285_297# VDD 3.2e-32
C128 sky130_fd_sc_hd__xor2_1_0/a_117_297# SUB -0.00177f
C129 VDD G3 0.0413f
C130 G3 G2 -1.94e-25
C131 A4 sky130_fd_sc_hd__and2_1_3/a_59_75# 0.0591f
C132 VDD sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.00867f
C133 sky130_fd_sc_hd__xor2_1_1/a_285_47# B2 2.25e-19
C134 sky130_fd_sc_hd__xor2_1_0/a_35_297# B1 0.0359f
C135 sky130_fd_sc_hd__xor2_1_3/a_35_297# A4 0.0402f
C136 sky130_fd_sc_hd__xor2_1_0/a_35_297# G2 2.05e-19
C137 sky130_fd_sc_hd__xor2_1_2/a_285_297# P2 2.5e-20
C138 B3 A4 0.00861f
C139 A2 A3 0.00809f
C140 P2 A3 0.00732f
C141 VDD sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.00949f
C142 G3 sky130_fd_sc_hd__and2_1_3/a_59_75# 9.08e-20
C143 VDD sky130_fd_sc_hd__xor2_1_3/a_117_297# -1.39e-19
C144 sky130_fd_sc_hd__xor2_1_1/a_35_297# G2 0.0663f
C145 sky130_fd_sc_hd__xor2_1_0/a_117_297# VDD -1.39e-19
C146 G3 sky130_fd_sc_hd__xor2_1_3/a_35_297# 5.99e-22
C147 A4 B4 0.249f
C148 B3 G3 0.0409f
C149 sky130_fd_sc_hd__xor2_1_0/a_117_297# G2 1.14e-19
C150 A4 sky130_fd_sc_hd__xor2_1_2/a_35_297# 0.0101f
C151 B2 sky130_fd_sc_hd__and2_1_0/a_59_75# 5.54e-20
C152 sky130_fd_sc_hd__xor2_1_2/a_117_297# SUB -0.00177f
C153 sky130_fd_sc_hd__xor2_1_3/a_285_297# B4 1.19e-19
C154 P1 sky130_fd_sc_hd__xor2_1_1/a_117_297# 1.21e-19
C155 G3 B4 3.51e-20
C156 sky130_fd_sc_hd__and2_1_1/a_59_75# B2 0.0564f
C157 G3 sky130_fd_sc_hd__xor2_1_2/a_35_297# 0.0665f
C158 B3 sky130_fd_sc_hd__xor2_1_1/a_35_297# 4e-19
C159 sky130_fd_sc_hd__and2_1_2/a_145_75# VDD -6.31e-19
C160 VDD sky130_fd_sc_hd__xor2_1_2/a_117_297# -1.39e-19
C161 P3 P4 2.91e-20
C162 SUB sky130_fd_sc_hd__xor2_1_1/a_117_297# -0.00177f
C163 P1 sky130_fd_sc_hd__xor2_1_1/a_285_297# 1.46e-19
C164 B2 sky130_fd_sc_hd__xor2_1_0/a_285_47# 5.6e-20
C165 P1 G1 3.4e-19
C166 B2 A3 0.00246f
C167 G3 P2 0.00384f
C168 B3 sky130_fd_sc_hd__and2_1_2/a_145_75# 2.46e-20
C169 VDD sky130_fd_sc_hd__and2_1_0/a_145_75# -6.31e-19
C170 A2 sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.0101f
C171 sky130_fd_sc_hd__xor2_1_0/a_35_297# P2 2.9e-21
C172 P1 SUB 0.0117f
C173 sky130_fd_sc_hd__and2_1_1/a_59_75# A3 3.22e-20
C174 sky130_fd_sc_hd__xor2_1_2/a_285_297# P4 2.02e-20
C175 A3 P4 3.19e-21
C176 sky130_fd_sc_hd__xor2_1_2/a_285_297# P3 0.00179f
C177 A2 sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.0397f
C178 VDD sky130_fd_sc_hd__xor2_1_1/a_117_297# -1.39e-19
C179 sky130_fd_sc_hd__xor2_1_1/a_35_297# P2 0.00234f
C180 A3 P3 0.006f
C181 sky130_fd_sc_hd__and2_1_2/a_59_75# SUB 0.00617f
C182 G2 sky130_fd_sc_hd__xor2_1_1/a_117_297# 7.26e-19
C183 G4 P4 0.00346f
C184 G1 SUB 0.00116f
C185 P3 G4 5.33e-19
C186 A1 sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.0402f
C187 VDD P1 0.0465f
C188 P1 B1 0.0021f
C189 P1 G2 6.62e-19
C190 VDD sky130_fd_sc_hd__and2_1_2/a_59_75# 0.00479f
C191 sky130_fd_sc_hd__xor2_1_2/a_285_297# A3 6.24e-19
C192 sky130_fd_sc_hd__xor2_1_0/a_117_297# A1 0.00414f
C193 VDD sky130_fd_sc_hd__xor2_1_1/a_285_297# 6.02e-20
C194 VDD G1 0.0385f
C195 B1 G1 0.0397f
C196 sky130_fd_sc_hd__xor2_1_2/a_285_297# G4 3.71e-19
C197 G2 sky130_fd_sc_hd__xor2_1_1/a_285_297# 5.75e-19
C198 A3 G4 1.26e-19
C199 G2 G1 0.00179f
C200 sky130_fd_sc_hd__xor2_1_2/a_117_297# P2 1.97e-20
C201 A4 P4 0.00232f
C202 A4 P3 0.0296f
C203 VDD SUB -0.222f
C204 B2 sky130_fd_sc_hd__xor2_1_0/a_35_297# 7.19e-19
C205 B1 SUB 0.134f
C206 B3 sky130_fd_sc_hd__and2_1_2/a_59_75# 0.0565f
C207 VDD sky130_fd_sc_hd__and2_1_1/a_145_75# -6.31e-19
C208 G2 SUB -1.95e-19
C209 sky130_fd_sc_hd__xor2_1_0/a_35_297# sky130_fd_sc_hd__and2_1_0/a_59_75# 5.6e-19
C210 sky130_fd_sc_hd__xor2_1_3/a_285_297# P4 0.0109f
C211 B2 sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.0446f
C212 sky130_fd_sc_hd__xor2_1_3/a_285_297# P3 9.07e-20
C213 G3 P3 2.77e-19
C214 sky130_fd_sc_hd__and2_1_1/a_59_75# sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.00179f
C215 sky130_fd_sc_hd__and2_1_3/a_59_75# SUB 0.00649f
C216 sky130_fd_sc_hd__xor2_1_2/a_35_297# sky130_fd_sc_hd__and2_1_2/a_59_75# 5.6e-19
C217 VDD sky130_fd_sc_hd__and2_1_3/a_145_75# -6.31e-19
C218 sky130_fd_sc_hd__xor2_1_3/a_35_297# SUB -0.0066f
C219 sky130_fd_sc_hd__xor2_1_2/a_285_297# A4 3.31e-19
C220 sky130_fd_sc_hd__and2_1_1/a_59_75# sky130_fd_sc_hd__xor2_1_1/a_35_297# 5.6e-19
C221 VDD B1 0.00679f
C222 A2 sky130_fd_sc_hd__xor2_1_1/a_117_297# 0.00414f
C223 A4 A3 0.00249f
C224 P2 sky130_fd_sc_hd__xor2_1_1/a_117_297# 5.63e-19
C225 B3 SUB 0.232f
C226 sky130_fd_sc_hd__xor2_1_1/a_35_297# P3 1.16e-20
C227 VDD G2 0.0388f
C228 sky130_fd_sc_hd__xor2_1_3/a_117_297# P4 5.63e-19
C229 B1 G2 8.95e-20
C230 sky130_fd_sc_hd__xor2_1_3/a_117_297# P3 7.54e-20
C231 sky130_fd_sc_hd__xor2_1_2/a_285_297# G3 6.58e-19
C232 A4 G4 0.0729f
C233 B4 SUB 0.154f
C234 A1 sky130_fd_sc_hd__and2_1_0/a_145_75# 0.00119f
C235 G3 A3 0.074f
C236 VDD sky130_fd_sc_hd__and2_1_3/a_59_75# -7.45e-19
C237 A2 P1 0.0305f
C238 sky130_fd_sc_hd__and2_1_2/a_145_75# B2 2.37e-21
C239 P1 P2 3.79e-19
C240 sky130_fd_sc_hd__xor2_1_2/a_35_297# SUB -0.0109f
C241 VDD sky130_fd_sc_hd__xor2_1_3/a_35_297# 0.00289f
C242 B3 sky130_fd_sc_hd__and2_1_3/a_145_75# 6.15e-21
C243 sky130_fd_sc_hd__xor2_1_3/a_285_297# G4 6.56e-19
C244 G3 G4 0.00197f
C245 B3 VDD 0.0264f
C246 P2 sky130_fd_sc_hd__and2_1_2/a_59_75# 0.00164f
C247 sky130_fd_sc_hd__xor2_1_1/a_35_297# A3 0.00595f
C248 B4 sky130_fd_sc_hd__and2_1_3/a_145_75# 2.46e-20
C249 A2 sky130_fd_sc_hd__xor2_1_1/a_285_297# 6.41e-19
C250 P2 sky130_fd_sc_hd__xor2_1_1/a_285_297# 0.0109f
C251 VDD B4 0.00646f
C252 A2 G1 1.33e-19
C253 A1 P1 0.00719f
C254 sky130_fd_sc_hd__xor2_1_3/a_35_297# sky130_fd_sc_hd__and2_1_3/a_59_75# 5.6e-19
C255 VDD sky130_fd_sc_hd__xor2_1_2/a_35_297# 0.0079f
C256 sky130_fd_sc_hd__xor2_1_0/a_285_297# P1 0.00448f
C257 G1 0 0.0305f
C258 SUB 0 2.81f
C259 VDD 0 7.09f
C260 P3 0 0.0173f
C261 sky130_fd_sc_hd__xor2_1_2/a_285_297# 0 0.00137f
C262 sky130_fd_sc_hd__xor2_1_2/a_35_297# 0 0.255f
C263 P2 0 0.0182f
C264 A2 0 0.317f
C265 B2 0 0.338f
C266 sky130_fd_sc_hd__xor2_1_1/a_285_297# 0 0.00137f
C267 sky130_fd_sc_hd__xor2_1_1/a_35_297# 0 0.255f
C268 P1 0 0.0183f
C269 A1 0 0.373f
C270 B1 0 0.337f
C271 sky130_fd_sc_hd__xor2_1_0/a_285_297# 0 0.00137f
C272 sky130_fd_sc_hd__xor2_1_0/a_35_297# 0 0.255f
C273 G4 0 0.0255f
C274 B4 0 0.342f
C275 A4 0 0.328f
C276 sky130_fd_sc_hd__and2_1_3/a_59_75# 0 0.177f
C277 G3 0 0.0256f
C278 B3 0 0.339f
C279 A3 0 0.323f
C280 sky130_fd_sc_hd__and2_1_2/a_59_75# 0 0.177f
C281 G2 0 0.0255f
C282 sky130_fd_sc_hd__and2_1_1/a_59_75# 0 0.177f
C283 sky130_fd_sc_hd__and2_1_0/a_59_75# 0 0.177f
C284 P4 0 0.0763f
C285 sky130_fd_sc_hd__xor2_1_3/a_285_297# 0 0.00137f
C286 sky130_fd_sc_hd__xor2_1_3/a_35_297# 0 0.255f
.ends

.subckt adder_4 A1 B1 A2 B2 S1 S2 S3 S4 CO VDD adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75#
+ adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_384_47# adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# adder_2_0/sky130_fd_sc_hd__a21o_1_2/X
+ adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_47#
+ adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75#
+ adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297#
+ adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_384_47#
+ adder_2_0/sky130_fd_sc_hd__and4_1_0/X adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297#
+ adder_3_0/G3 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# adder_3_0/G2 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B
+ adder_3_0/G1 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297#
+ adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_3_0/sky130_fd_sc_hd__xor2_1_1/B
+ adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21#
+ A4 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_47# A3 adder_3_0/P4 B4 B3 adder_1_0/sky130_fd_sc_hd__and2_1_3/a_145_75#
+ adder_3_0/P3 adder_3_0/P2 CI adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# adder_3_0/P1
+ adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297#
+ SUB adder_2_0/G4
Xadder_2_0 CI adder_3_0/P1 adder_3_0/G1 adder_3_0/P2 adder_3_0/G2 adder_3_0/P3 adder_3_0/G3
+ adder_3_0/P4 adder_2_0/G4 CO adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47#
+ adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_384_47# adder_2_0/sky130_fd_sc_hd__a21o_1_1/X
+ adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21#
+ VDD adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_384_47#
+ adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# adder_2_0/sky130_fd_sc_hd__and4_1_0/a_109_47#
+ adder_2_0/sky130_fd_sc_hd__a21o_1_2/X adder_2_0/sky130_fd_sc_hd__a21o_1_0/X adder_2_0/sky130_fd_sc_hd__and4_1_0/X
+ adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21#
+ SUB adder_2_0/sky130_fd_sc_hd__and4_1_0/a_197_47# adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_384_47#
+ adder_2_0/sky130_fd_sc_hd__and4_1_0/a_303_47# adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21#
+ adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_384_47# adder_2
Xadder_3_0 adder_3_0/G1 adder_3_0/P2 adder_3_0/G2 adder_3_0/G3 adder_3_0/P4 S1 S2
+ S3 S4 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_117_297# adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297#
+ adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_47#
+ adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_384_47#
+ adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297#
+ adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_47# adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_299_297#
+ adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297#
+ adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297#
+ adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297#
+ adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_47#
+ adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21#
+ adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_384_47# adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_117_297#
+ adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_47#
+ adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_117_297# CI adder_3_0/P1 SUB adder_3_0/sky130_fd_sc_hd__xor2_1_2/B
+ adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# VDD adder_3_0/P3 adder_3
Xadder_1_0 A1 B1 A2 B2 A3 B3 A4 B4 adder_3_0/G1 adder_3_0/P1 adder_3_0/G2 adder_3_0/P2
+ adder_3_0/G3 adder_3_0/P3 adder_2_0/G4 adder_3_0/P4 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_117_297#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_47#
+ adder_1_0/sky130_fd_sc_hd__and2_1_3/a_145_75# adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_47#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# adder_1_0/sky130_fd_sc_hd__and2_1_0/a_145_75#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_47#
+ adder_1_0/sky130_fd_sc_hd__and2_1_1/a_145_75# adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_47# adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_117_297#
+ adder_1_0/sky130_fd_sc_hd__and2_1_2/a_145_75# SUB adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# VDD adder_1
C0 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# 1.09e-19
C1 adder_3_0/P3 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.00106f
C2 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# adder_3_0/P1 0.0174f
C3 SUB B2 0.00396f
C4 CO adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# 4.34e-19
C5 VDD adder_3_0/G2 0.293f
C6 A3 B1 9.01e-19
C7 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_3_0/sky130_fd_sc_hd__xor2_1_2/B -0.00531f
C8 B3 B1 5.26e-19
C9 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# CI 3.01e-20
C10 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# adder_3_0/P3 -0.00186f
C11 adder_3_0/G1 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 0.0407f
C12 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# adder_3_0/G2 7.19e-20
C13 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# adder_3_0/P3 0.00147f
C14 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 6.98e-20
C15 SUB adder_3_0/sky130_fd_sc_hd__xor2_1_2/B -0.00596f
C16 S1 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 5.99e-19
C17 adder_2_0/G4 adder_3_0/P1 0.03f
C18 adder_2_0/sky130_fd_sc_hd__and4_1_0/X adder_2_0/sky130_fd_sc_hd__a21o_1_2/X -0.0153f
C19 adder_3_0/P3 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 0.00405f
C20 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# adder_3_0/sky130_fd_sc_hd__xor2_1_2/B -0.00349f
C21 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X A1 2.52e-21
C22 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_3_0/G3 0.0147f
C23 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# A4 -2.86e-19
C24 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# adder_3_0/G3 1.82e-20
C25 S4 S1 0.0283f
C26 adder_3_0/P2 CI 0.0316f
C27 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_3_0/G2 1.77e-21
C28 adder_3_0/G1 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.00976f
C29 B4 adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 5.56e-19
C30 adder_2_0/G4 A3 2.73e-19
C31 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_3_0/P2 0.00226f
C32 adder_3_0/G2 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 2.92e-19
C33 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_384_47# CI 1.5e-20
C34 adder_2_0/G4 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 1.23e-20
C35 adder_3_0/P1 A3 1.31e-19
C36 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 2.84e-20
C37 adder_2_0/G4 B3 2.86e-19
C38 adder_3_0/P3 adder_3_0/G3 0.318f
C39 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# CI 0.00104f
C40 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# B2 6.16e-19
C41 adder_3_0/P1 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# -9.58e-19
C42 A2 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.00125f
C43 adder_3_0/P4 adder_3_0/P2 0.0172f
C44 adder_1_0/sky130_fd_sc_hd__and2_1_3/a_145_75# adder_3_0/P3 6.88e-19
C45 B3 adder_3_0/P1 1.06e-19
C46 S3 S2 0.717f
C47 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X SUB 6.92e-20
C48 adder_3_0/G2 adder_3_0/P3 0.0027f
C49 A4 CI 0.0346f
C50 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 2.6e-20
C51 adder_3_0/P4 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_47# 5.65e-19
C52 SUB adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 3.16e-20
C53 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# adder_3_0/sky130_fd_sc_hd__xor2_1_1/B -3.51e-21
C54 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 6.84e-21
C55 B3 A3 1.3f
C56 adder_3_0/P2 B2 0.0325f
C57 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_3_0/sky130_fd_sc_hd__xor2_1_3/B -0.00152f
C58 adder_3_0/G1 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 3.22e-19
C59 adder_3_0/P4 A4 0.00541f
C60 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# adder_3_0/P2 2.5e-19
C61 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_47# adder_3_0/P2 0.00105f
C62 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 1.13e-19
C63 adder_3_0/G1 B4 6.45e-20
C64 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_384_47# CI 6.1e-19
C65 A2 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0.00352f
C66 S2 SUB 0.089f
C67 VDD A1 0.37f
C68 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_3_0/P2 -0.0409f
C69 B4 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 3.05e-20
C70 CO adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.00229f
C71 A4 B2 8.41e-19
C72 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# SUB -5.69e-20
C73 A2 B4 3.27e-19
C74 VDD adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 3.54e-19
C75 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_3_0/G3 0.0318f
C76 S4 CO 0.209f
C77 adder_2_0/G4 adder_2_0/sky130_fd_sc_hd__and4_1_0/X 1.36e-19
C78 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_3_0/G2 0.0309f
C79 VDD S4 -2.22e-19
C80 adder_2_0/sky130_fd_sc_hd__and4_1_0/X adder_3_0/P1 0.00468f
C81 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# B4 3.05e-20
C82 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# B1 3.89e-20
C83 S1 CO 0.257f
C84 VDD adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 6.51e-19
C85 adder_3_0/G1 SUB 0.376f
C86 adder_2_0/G4 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 1.9e-19
C87 VDD S1 -0.00144f
C88 B4 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 5.38e-20
C89 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_3_0/G3 0.00129f
C90 SUB adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 3.52e-21
C91 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 8.63e-21
C92 adder_3_0/P3 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 4.09e-20
C93 S3 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# -7.21e-19
C94 adder_2_0/sky130_fd_sc_hd__and4_1_0/X A3 3.53e-20
C95 adder_3_0/P2 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 1.63e-19
C96 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X CI 0.0104f
C97 A2 SUB 0.00582f
C98 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X adder_3_0/P2 0.00437f
C99 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_3_0/G2 0.00105f
C100 adder_2_0/sky130_fd_sc_hd__and4_1_0/X adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 1.35e-19
C101 S3 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 0.00612f
C102 VDD adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 0.00147f
C103 B3 adder_2_0/sky130_fd_sc_hd__and4_1_0/X 1.55e-20
C104 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# A3 -7.46e-20
C105 adder_2_0/G4 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# 5.98e-20
C106 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# SUB 1.84e-20
C107 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_117_297# adder_3_0/G3 -9e-22
C108 B3 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 0.0107f
C109 adder_3_0/P4 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 0.0226f
C110 adder_2_0/G4 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 0.00256f
C111 SUB adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# -2.23e-19
C112 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# S1 -1.76e-19
C113 adder_3_0/P4 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 0.00101f
C114 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_3_0/P1 0.00383f
C115 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_3_0/P3 0.00801f
C116 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_3_0/P1 -6.47e-19
C117 B3 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_47# 5.14e-19
C118 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# adder_3_0/G3 3.83e-19
C119 SUB adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 8.85e-19
C120 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# adder_3_0/G3 0.00128f
C121 S2 adder_3_0/P2 0.0771f
C122 B2 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 1.92e-20
C123 adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# A4 0.0161f
C124 S4 adder_3_0/P3 -8.8e-19
C125 adder_3_0/G1 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 3.92e-20
C126 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 9.58e-21
C127 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# SUB 0.00127f
C128 B3 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# 0.00199f
C129 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# adder_3_0/G2 1.95e-19
C130 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_3_0/P3 5.63e-21
C131 B4 adder_3_0/G3 9.64e-20
C132 S1 adder_3_0/P3 0.1f
C133 SUB adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# -5.95e-20
C134 B1 CI 1.95e-19
C135 A2 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 0.0155f
C136 B4 adder_3_0/G2 9.64e-20
C137 adder_2_0/G4 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 0.00895f
C138 adder_3_0/P4 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_47# 0.00104f
C139 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# CI 0.00244f
C140 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 4.82e-20
C141 adder_3_0/G1 adder_3_0/P2 0.268f
C142 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X adder_3_0/P3 0.024f
C143 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_3_0/G3 0.00131f
C144 VDD CO 0.114f
C145 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 2.84e-32
C146 adder_3_0/G1 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_384_47# 1.56e-20
C147 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_47# adder_3_0/sky130_fd_sc_hd__xor2_1_2/B -5.8e-19
C148 adder_3_0/P2 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 0.00223f
C149 adder_2_0/G4 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 9.53e-20
C150 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_3_0/G2 0.0146f
C151 A2 adder_3_0/P2 0.00581f
C152 SUB adder_3_0/G3 1.22f
C153 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_3_0/G1 0.0239f
C154 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# adder_3_0/P4 -2.26e-19
C155 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# adder_3_0/G3 4.76e-20
C156 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# -9.51e-19
C157 S1 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# -3.09e-20
C158 SUB adder_3_0/G2 0.287f
C159 adder_2_0/G4 CI 0.0329f
C160 adder_3_0/G1 A4 7.97e-20
C161 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# adder_3_0/G2 0.00591f
C162 B1 B2 0.00145f
C163 adder_2_0/G4 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.00465f
C164 adder_3_0/P1 CI 0.154f
C165 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# A1 -6.08e-19
C166 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 6.41e-20
C167 A4 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 3.72e-20
C168 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_3_0/P1 5.66e-20
C169 adder_3_0/P2 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.0148f
C170 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# B2 5.71e-20
C171 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# adder_3_0/G3 0.00552f
C172 A2 A4 4.9e-19
C173 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B S1 0.00968f
C174 adder_3_0/G1 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_47# 6.94e-19
C175 adder_2_0/G4 adder_3_0/P4 1.29f
C176 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 6.98e-20
C177 VDD adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 1.34e-19
C178 A3 CI 0.0954f
C179 adder_3_0/P4 adder_3_0/P1 0.0308f
C180 VDD adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 5.68e-32
C181 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# CI 0.00503f
C182 adder_2_0/sky130_fd_sc_hd__and4_1_0/X adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 6.46e-21
C183 B3 CI 0.208f
C184 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# A4 3.72e-20
C185 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 5.75e-20
C186 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 2.45e-19
C187 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 2.82e-21
C188 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_384_47# adder_3_0/P1 5.17e-19
C189 CO adder_3_0/P3 0.0888f
C190 adder_2_0/G4 B2 0.00161f
C191 A4 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 6.49e-20
C192 B4 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 0.0072f
C193 adder_3_0/P2 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# -1.11e-20
C194 adder_3_0/P4 A3 1.54e-19
C195 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_3_0/G3 0.00261f
C196 VDD adder_3_0/P3 0.534f
C197 adder_3_0/P1 B2 0.00166f
C198 adder_3_0/P4 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 1.49e-19
C199 B3 adder_3_0/P4 1.46e-19
C200 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_3_0/G2 0.0173f
C201 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 5.31e-21
C202 S2 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 0.00273f
C203 S2 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_47# 9.42e-19
C204 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_145_75# adder_3_0/G3 1.86e-19
C205 B4 A1 2.13e-19
C206 A3 B2 0.938f
C207 adder_2_0/G4 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 8.62e-20
C208 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X B1 2.31e-20
C209 adder_3_0/P2 adder_3_0/G3 0.771f
C210 A4 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 0.00264f
C211 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_3_0/P1 0.103f
C212 adder_3_0/G2 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_145_75# 8.25e-19
C213 B3 B2 0.00119f
C214 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 1.53e-19
C215 CO adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 6.62e-19
C216 adder_3_0/G1 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 3.53e-20
C217 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# adder_3_0/P3 1.5e-20
C218 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_384_47# 7.63e-20
C219 adder_3_0/P2 adder_3_0/G2 0.749f
C220 S3 S4 0.442f
C221 S1 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# 1.21e-20
C222 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_3_0/P3 0.00509f
C223 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_384_47# 7.89e-20
C224 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 8.48e-19
C225 adder_3_0/P3 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 1.27e-21
C226 S3 S1 0.0279f
C227 A2 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 2.61e-19
C228 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# -0.00268f
C229 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_3_0/G2 0.00723f
C230 SUB A1 0.00365f
C231 adder_2_0/sky130_fd_sc_hd__and4_1_0/X CI 0.0231f
C232 A4 adder_3_0/G3 1.67e-19
C233 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B CO 0.0577f
C234 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_117_297# S1 -4.4e-19
C235 VDD adder_3_0/sky130_fd_sc_hd__xor2_1_1/B -0.0577f
C236 A4 adder_3_0/G2 1.16e-19
C237 SUB adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 7.61e-19
C238 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# CI 0.0185f
C239 adder_3_0/P1 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 5.1e-19
C240 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X adder_3_0/P1 0.0283f
C241 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_47# adder_3_0/G3 0.00103f
C242 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_117_297# adder_3_0/P2 0.00103f
C243 adder_2_0/G4 adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 0.0161f
C244 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 3.35e-21
C245 adder_3_0/P4 adder_2_0/sky130_fd_sc_hd__and4_1_0/X 2.22e-19
C246 S4 SUB 0.0982f
C247 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_47# CI 9.49e-19
C248 S4 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_117_297# -3.24e-19
C249 SUB adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 4.5e-19
C250 adder_3_0/P1 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_197_47# 2.07e-19
C251 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_3_0/P4 5.92e-20
C252 SUB S1 1.14f
C253 VDD adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# -4.41e-19
C254 adder_3_0/G1 B1 0.087f
C255 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 9.14e-21
C256 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# S1 -6.35e-20
C257 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# CI 0.00225f
C258 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# -8.36e-21
C259 adder_2_0/G4 S2 2.28e-20
C260 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# CI 2.82e-19
C261 adder_3_0/P3 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 3.13e-19
C262 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B CI 1.31e-19
C263 SUB adder_2_0/sky130_fd_sc_hd__a21o_1_1/X -6.74e-19
C264 A2 B1 0.403f
C265 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 7.55e-22
C266 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_303_47# CO 5.64e-19
C267 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# adder_3_0/P1 0.00143f
C268 CO adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# 0.00874f
C269 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# B1 6.38e-19
C270 adder_2_0/sky130_fd_sc_hd__and4_1_0/X adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 6.99e-21
C271 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_3_0/P3 0.131f
C272 adder_3_0/P4 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 0.0108f
C273 VDD adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# 0.00215f
C274 adder_2_0/G4 adder_3_0/G1 3.67e-20
C275 S3 CO 0.119f
C276 VDD adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 5.68e-32
C277 S2 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.00567f
C278 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X adder_3_0/G3 0.0333f
C279 adder_3_0/G1 adder_3_0/P1 0.0488f
C280 A1 adder_3_0/P2 3.75e-19
C281 S3 VDD 8.27e-19
C282 adder_2_0/G4 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 4.89e-20
C283 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 4.7e-20
C284 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_117_297# CO 0.00216f
C285 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 1.5e-20
C286 adder_3_0/G2 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 1.74e-19
C287 B3 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# 4.93e-21
C288 VDD B4 0.138f
C289 adder_2_0/G4 A2 1.33e-19
C290 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_3_0/P2 -8.11e-19
C291 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_3_0/P3 5.23e-19
C292 A2 adder_3_0/P1 0.0449f
C293 adder_3_0/G1 A3 1.32e-19
C294 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# A1 9.74e-19
C295 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_145_75# adder_3_0/G3 8.23e-19
C296 adder_3_0/P4 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 0.0131f
C297 B3 adder_3_0/G1 1.01e-19
C298 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 4.59e-19
C299 A3 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 0.0163f
C300 VDD adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 6.69e-20
C301 A1 A4 2.8e-19
C302 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# adder_3_0/P1 -6e-21
C303 A2 A3 0.00214f
C304 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 3.66e-20
C305 adder_2_0/G4 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 7.97e-20
C306 S1 adder_3_0/P2 0.234f
C307 S4 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_47# 0.00104f
C308 SUB CO 0.151f
C309 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_3_0/sky130_fd_sc_hd__xor2_1_2/B -0.0029f
C310 B3 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 4.89e-20
C311 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_117_297# adder_3_0/P3 3.36e-20
C312 adder_3_0/P1 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 1.38e-19
C313 VDD SUB 1.2f
C314 B3 A2 7.94e-19
C315 adder_3_0/P4 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 5.12e-19
C316 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# CI 2.83e-19
C317 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 0.00309f
C318 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_303_47# adder_3_0/P3 4e-19
C319 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# A3 5.96e-20
C320 adder_2_0/sky130_fd_sc_hd__and4_1_0/X adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 5.71e-20
C321 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X adder_3_0/P2 0.0193f
C322 adder_2_0/G4 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 1.03e-19
C323 B1 adder_3_0/G3 0.00439f
C324 adder_2_0/G4 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 0.00559f
C325 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# adder_3_0/P3 1.34e-19
C326 A3 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 5.49e-19
C327 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# B3 4.65e-20
C328 adder_3_0/P4 CI 0.0664f
C329 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# adder_3_0/G3 3.99e-20
C330 adder_3_0/G2 B1 0.00409f
C331 adder_2_0/G4 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 1.65e-19
C332 S3 adder_3_0/P3 0.0899f
C333 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_3_0/P4 4.73e-19
C334 S2 adder_2_0/sky130_fd_sc_hd__and4_1_0/X 1.66e-20
C335 B3 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 2.25e-20
C336 B4 adder_3_0/P3 0.00132f
C337 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_384_47# CI 2.66e-19
C338 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_117_297# adder_3_0/P3 1.69e-19
C339 SUB adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 4.59e-19
C340 B2 CI 3.41e-19
C341 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# B2 8.1e-20
C342 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# adder_3_0/P2 0.00724f
C343 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# -7.49e-19
C344 adder_2_0/G4 adder_3_0/G3 0.217f
C345 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_3_0/P3 1.7e-19
C346 B3 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 0.0195f
C347 adder_2_0/G4 adder_1_0/sky130_fd_sc_hd__and2_1_3/a_145_75# 8.23e-19
C348 adder_3_0/P1 adder_3_0/G3 0.197f
C349 VDD adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 2.99e-19
C350 adder_3_0/P4 B2 6.88e-19
C351 adder_2_0/G4 adder_3_0/G2 7.19e-19
C352 adder_2_0/sky130_fd_sc_hd__and4_1_0/X adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 7.41e-22
C353 SUB adder_3_0/P3 0.136f
C354 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B CI -0.005f
C355 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_384_47# adder_3_0/P2 4.8e-19
C356 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_384_47# adder_3_0/G3 4.39e-19
C357 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# adder_3_0/P3 0.00176f
C358 adder_3_0/P1 adder_3_0/G2 0.405f
C359 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 4.77e-19
C360 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# 0.00254f
C361 A3 adder_3_0/G3 0.0807f
C362 S2 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 0.0283f
C363 adder_3_0/G2 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_384_47# 7.32e-20
C364 CO adder_3_0/P2 0.108f
C365 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 9.34e-21
C366 S3 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B -1.33e-20
C367 VDD adder_3_0/P2 0.267f
C368 A3 adder_3_0/G2 2.08e-19
C369 B3 adder_3_0/G3 0.0363f
C370 adder_3_0/P4 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 4.82e-19
C371 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# adder_3_0/P3 0.0105f
C372 B3 adder_3_0/G2 1.49e-19
C373 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_47# adder_3_0/P3 1.14e-19
C374 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# VDD 0.00637f
C375 S1 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 6.31e-20
C376 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_117_297# adder_3_0/P1 3.02e-21
C377 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X CI 0.00101f
C378 S1 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 3.79e-19
C379 VDD A4 0.142f
C380 B4 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 5.38e-20
C381 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# adder_3_0/sky130_fd_sc_hd__xor2_1_2/B -2.17e-19
C382 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# adder_3_0/P2 0.00132f
C383 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_3_0/P2 0.00106f
C384 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_3_0/P3 5.59e-20
C385 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_117_297# A3 2.11e-19
C386 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B SUB 0.00204f
C387 A1 B1 0.237f
C388 adder_3_0/P2 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 0.0124f
C389 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# CI 0.00313f
C390 CO adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_384_47# 3.28e-19
C391 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_117_297# B4 0.00366f
C392 adder_2_0/G4 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 2.44e-19
C393 adder_3_0/P4 adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 4.95e-20
C394 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.00238f
C395 S2 CI 0.00387f
C396 adder_3_0/P2 adder_3_0/P3 0.405f
C397 SUB adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# -5.32e-19
C398 adder_3_0/P4 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 4.86e-19
C399 adder_2_0/sky130_fd_sc_hd__and4_1_0/X adder_3_0/G3 4.68e-20
C400 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 2.85e-19
C401 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# CI 0.0208f
C402 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_47# adder_3_0/P3 -3.53e-19
C403 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_109_47# CI 3.82e-20
C404 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_3_0/G3 0.00202f
C405 S2 adder_3_0/P4 9.76e-19
C406 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# S1 9.19e-19
C407 A1 adder_3_0/P1 0.00472f
C408 adder_2_0/G4 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 1.01e-20
C409 adder_3_0/G1 CI 0.0965f
C410 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X B1 3.97e-19
C411 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_3_0/G2 1.11e-21
C412 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 1.8e-19
C413 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# adder_3_0/P4 1.73e-19
C414 A4 adder_3_0/P3 0.0462f
C415 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 3.33e-20
C416 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_3_0/P1 7.47e-19
C417 CO adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 0.0284f
C418 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# CI 5.48e-19
C419 A1 A3 5.77e-19
C420 A2 CI 2.43e-19
C421 SUB adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# 1.4e-19
C422 VDD adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 0.00224f
C423 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# adder_3_0/G3 3.28e-19
C424 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# CO 7.73e-19
C425 adder_3_0/G1 adder_3_0/P4 1.36e-20
C426 B3 A1 3.87e-19
C427 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# A2 9.74e-19
C428 adder_2_0/G4 S1 2.86e-20
C429 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_3_0/P1 7.78e-20
C430 S3 SUB 0.0872f
C431 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_3_0/G3 0.00395f
C432 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_3_0/G3 0.0127f
C433 S1 adder_3_0/P1 0.0451f
C434 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# CI 2.96e-20
C435 adder_3_0/P4 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 3.55e-20
C436 SUB B4 0.00678f
C437 adder_3_0/G1 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_384_47# 4.44e-19
C438 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_3_0/P2 0.0337f
C439 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_3_0/G2 0.0185f
C440 A2 adder_3_0/P4 4.36e-19
C441 S2 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.118f
C442 adder_2_0/G4 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 0.0203f
C443 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# CI 4.53e-20
C444 adder_3_0/G1 B2 2.02e-19
C445 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X adder_3_0/P1 0.0208f
C446 SUB adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 4.55e-19
C447 S1 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# -0.00115f
C448 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 9.82e-21
C449 A2 B2 0.77f
C450 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_3_0/P2 2.17e-19
C451 S3 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_47# 9.42e-19
C452 adder_3_0/P4 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 7.7e-20
C453 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# adder_3_0/G3 -5.99e-22
C454 adder_3_0/G1 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B -6.76e-19
C455 CI adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 0.00281f
C456 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# adder_3_0/P4 0.0141f
C457 VDD B1 0.244f
C458 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# B2 7.88e-20
C459 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# CO 0.00806f
C460 adder_3_0/P3 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 0.0225f
C461 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# adder_3_0/P4 0.00776f
C462 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# B2 0.0195f
C463 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# adder_3_0/G3 0.00432f
C464 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# adder_3_0/P1 0.00281f
C465 adder_3_0/P4 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 0.0105f
C466 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# VDD 0.00235f
C467 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# A4 6.49e-20
C468 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_3_0/P3 2.95e-20
C469 B4 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 3.05e-20
C470 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# B1 0.00429f
C471 adder_3_0/P4 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# -2.02e-20
C472 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_303_47# adder_3_0/P2 1.69e-19
C473 adder_3_0/G2 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 3.05e-20
C474 CI adder_3_0/G3 0.164f
C475 adder_3_0/P2 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# 0.00114f
C476 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# adder_3_0/P2 -1.01e-20
C477 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_3_0/G3 0.0177f
C478 adder_2_0/G4 CO 1.56e-19
C479 S3 adder_3_0/P2 3.05e-21
C480 adder_3_0/G2 CI 0.0259f
C481 adder_3_0/G1 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 0.0445f
C482 CO adder_3_0/P1 0.0294f
C483 adder_2_0/G4 VDD 0.174f
C484 B4 adder_3_0/P2 9.02e-20
C485 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_3_0/G2 9.85e-20
C486 S3 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_47# 7.3e-19
C487 adder_3_0/P4 adder_3_0/G3 0.00126f
C488 VDD adder_3_0/P1 0.332f
C489 SUB adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 1.84e-20
C490 S1 adder_2_0/sky130_fd_sc_hd__and4_1_0/X 0.00171f
C491 adder_3_0/P4 adder_3_0/G2 4.99e-20
C492 CO A3 0.00124f
C493 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 2.93e-19
C494 CO adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.014f
C495 adder_3_0/P4 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# 4.5e-19
C496 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# adder_3_0/P1 3.41e-19
C497 VDD A3 0.208f
C498 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_3_0/P2 0.00225f
C499 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# A1 0.00131f
C500 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 1.11e-19
C501 B2 adder_3_0/G3 0.00108f
C502 VDD adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 4.68e-19
C503 B4 A4 1.95f
C504 B3 VDD 0.171f
C505 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# adder_3_0/P3 0.00835f
C506 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# -4.45e-20
C507 SUB adder_3_0/P2 0.0707f
C508 adder_2_0/G4 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.00122f
C509 adder_3_0/G2 B2 0.089f
C510 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# adder_3_0/P1 0.00658f
C511 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# adder_3_0/P2 0.00898f
C512 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_3_0/P1 2.37e-21
C513 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_47# adder_3_0/G2 6.94e-19
C514 S4 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 0.00146f
C515 adder_3_0/P1 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 3.68e-21
C516 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# SUB 9.07e-20
C517 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_3_0/G3 0.00104f
C518 adder_3_0/G1 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_145_75# 0.00101f
C519 S1 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 0.0151f
C520 adder_2_0/G4 adder_3_0/P3 1.15f
C521 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_3_0/G2 0.0946f
C522 SUB A4 0.00516f
C523 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# adder_3_0/P2 0.00242f
C524 A3 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 9.09e-19
C525 adder_3_0/P1 adder_3_0/P3 0.649f
C526 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_2_0/sky130_fd_sc_hd__a21o_1_1/X -4.9e-21
C527 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_117_297# B2 0.00385f
C528 adder_3_0/P3 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_384_47# 4.84e-19
C529 adder_3_0/G1 A2 3.33e-19
C530 A3 adder_3_0/P3 0.002f
C531 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_3_0/P3 1.78e-19
C532 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 1.39e-20
C533 adder_3_0/P2 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 1.21e-19
C534 adder_3_0/P4 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 0.011f
C535 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X adder_3_0/G3 0.00133f
C536 CO adder_2_0/sky130_fd_sc_hd__and4_1_0/X 0.106f
C537 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# adder_3_0/G1 0.0212f
C538 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# S2 2.81e-19
C539 B3 adder_3_0/P3 0.0502f
C540 A1 CI 1.72e-19
C541 VDD adder_2_0/sky130_fd_sc_hd__and4_1_0/X -0.0032f
C542 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X adder_3_0/G2 0.0275f
C543 adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# adder_3_0/G3 2.97e-20
C544 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# CI 3.33e-19
C545 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# B1 0.022f
C546 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# A2 1.08e-19
C547 S3 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 0.00559f
C548 VDD adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# -6.68e-19
C549 S1 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# -2.34e-19
C550 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# adder_3_0/G3 1.39e-19
C551 A2 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 1.78e-19
C552 adder_2_0/G4 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 1.36e-19
C553 A4 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 3.72e-20
C554 VDD adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_47# -8.51e-21
C555 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# CI 0.0052f
C556 adder_3_0/P4 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 3.44e-19
C557 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_3_0/P1 0.0196f
C558 S1 CI 4.68e-19
C559 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 2.99e-20
C560 A1 B2 9.29e-19
C561 S4 adder_3_0/P4 0.0312f
C562 SUB adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 1.34e-19
C563 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# adder_3_0/G3 3.12e-19
C564 CO adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 0.0228f
C565 adder_3_0/P2 A4 1.08e-19
C566 VDD adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 0.00221f
C567 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X CI 2.11e-19
C568 VDD adder_3_0/sky130_fd_sc_hd__xor2_1_3/B -2.88e-19
C569 SUB adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 6.56e-19
C570 S1 adder_3_0/P4 0.00107f
C571 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# B1 0.00727f
C572 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_3_0/P1 0.0152f
C573 adder_3_0/G1 adder_3_0/G3 0.0163f
C574 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_145_75# adder_3_0/G2 5.09e-21
C575 adder_2_0/sky130_fd_sc_hd__and4_1_0/X adder_3_0/P3 5.85e-19
C576 B4 B1 2.5e-19
C577 adder_3_0/P4 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 0.00539f
C578 adder_2_0/G4 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_117_297# 3.36e-19
C579 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# A3 1e-19
C580 adder_3_0/G1 adder_3_0/G2 0.872f
C581 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_3_0/G3 0.0163f
C582 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_3_0/P3 0.011f
C583 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_3_0/sky130_fd_sc_hd__xor2_1_2/B -2.45e-19
C584 A2 adder_3_0/G3 0.0115f
C585 B3 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 7.98e-20
C586 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_3_0/G2 1.78e-20
C587 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# CI 4.51e-20
C588 A2 adder_3_0/G2 0.084f
C589 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_47# adder_3_0/P3 9.41e-19
C590 VDD adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# -9.12e-19
C591 S4 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.0035f
C592 adder_2_0/G4 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# 1.75e-19
C593 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X B2 2.07e-20
C594 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_3_0/sky130_fd_sc_hd__xor2_1_2/B -0.00197f
C595 adder_3_0/P1 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# 0.00112f
C596 S3 adder_2_0/G4 2.78e-20
C597 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# adder_3_0/P1 0.00383f
C598 S1 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.0236f
C599 CO adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 1.62e-20
C600 SUB B1 0.00716f
C601 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 2.6e-21
C602 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# adder_3_0/P3 1.03e-19
C603 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_3_0/G3 4.15e-19
C604 adder_2_0/G4 B4 0.0886f
C605 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# adder_3_0/G2 7.89e-19
C606 VDD adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# -0.00753f
C607 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X A1 2.97e-19
C608 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# SUB 1.54e-19
C609 B4 adder_3_0/P1 4.85e-20
C610 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_3_0/P3 5.91e-19
C611 A3 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# 2.34e-21
C612 adder_3_0/G2 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.00912f
C613 CO CI 0.0904f
C614 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_3_0/P3 -0.00685f
C615 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.00475f
C616 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 4.05e-20
C617 VDD CI 1.6f
C618 B3 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# 9.41e-19
C619 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_2_0/sky130_fd_sc_hd__and4_1_0/X 7.03e-19
C620 adder_3_0/P2 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 0.0208f
C621 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# VDD 0.00242f
C622 B4 A3 8.32e-19
C623 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# adder_3_0/G3 2.64e-19
C624 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_3_0/P1 5.85e-19
C625 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_3_0/P2 -4.84e-19
C626 adder_3_0/P4 CO 6.01e-19
C627 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 2.14e-20
C628 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# adder_3_0/G2 2.56e-19
C629 B3 B4 8.66e-19
C630 adder_2_0/G4 SUB 0.132f
C631 adder_2_0/G4 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_117_297# 3.67e-19
C632 VDD adder_3_0/P4 0.896f
C633 SUB adder_3_0/P1 0.175f
C634 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_145_75# adder_3_0/P2 4.99e-19
C635 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# adder_3_0/P1 1.85e-21
C636 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# adder_3_0/P3 3.07e-20
C637 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# CI 0.0137f
C638 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X adder_2_0/sky130_fd_sc_hd__a21o_1_1/X -9.62e-21
C639 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# CI 2.49e-19
C640 SUB A3 0.00693f
C641 VDD B2 0.176f
C642 S1 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# -7.29e-19
C643 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.0026f
C644 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# CO 8.7e-19
C645 SUB adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 8.68e-19
C646 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# adder_3_0/P3 0.0383f
C647 S2 S4 0.0289f
C648 adder_3_0/G2 adder_3_0/G3 0.882f
C649 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 3.16e-19
C650 B3 SUB 0.00596f
C651 adder_3_0/G1 A1 0.0955f
C652 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_3_0/sky130_fd_sc_hd__xor2_1_3/B -8.72e-21
C653 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# adder_3_0/P1 1.34e-20
C654 S2 S1 1.02f
C655 CO adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.477f
C656 adder_3_0/P2 B1 6.78e-19
C657 adder_3_0/P3 CI 0.132f
C658 adder_3_0/P4 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 2.19e-20
C659 VDD adder_3_0/sky130_fd_sc_hd__xor2_1_2/B -0.019f
C660 A2 A1 0.00288f
C661 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_3_0/P3 1.67e-19
C662 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# adder_3_0/P2 4.11e-19
C663 adder_2_0/G4 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 1.82e-19
C664 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 1.46e-20
C665 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# B1 8.1e-20
C666 adder_3_0/G1 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 0.017f
C667 adder_3_0/P1 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 0.00384f
C668 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# A1 0.0155f
C669 adder_3_0/P4 adder_3_0/P3 0.232f
C670 B2 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 0.00715f
C671 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_117_297# adder_3_0/G3 8.67e-21
C672 A4 B1 3.49e-19
C673 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# B4 -3.44e-20
C674 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_117_297# adder_3_0/G2 4.07e-19
C675 adder_2_0/G4 adder_3_0/P2 0.0231f
C676 A3 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 5.96e-20
C677 CO adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0.00661f
C678 adder_3_0/P1 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_145_75# 6.85e-19
C679 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# adder_3_0/sky130_fd_sc_hd__xor2_1_2/B -0.00512f
C680 adder_3_0/G1 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 1.03e-19
C681 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_3_0/sky130_fd_sc_hd__xor2_1_2/B -9.88e-19
C682 adder_3_0/P3 B2 0.00568f
C683 adder_3_0/P1 adder_3_0/P2 1.17f
C684 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# -0.00611f
C685 VDD adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# -5.68e-32
C686 VDD adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 0.0342f
C687 B3 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 4.65e-20
C688 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# adder_3_0/P3 0.00275f
C689 A2 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 1.47e-20
C690 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# 1.37e-21
C691 SUB adder_2_0/sky130_fd_sc_hd__and4_1_0/X 1.11e-19
C692 CO adder_2_0/sky130_fd_sc_hd__and4_1_0/a_197_47# 4.68e-19
C693 VDD adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# -5.1e-20
C694 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B CI 0.0245f
C695 adder_3_0/P4 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 0.00212f
C696 A3 adder_3_0/P2 0.0346f
C697 CO adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 0.00441f
C698 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_3_0/P1 0.00259f
C699 S4 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# -1.86e-19
C700 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_47# adder_3_0/P2 -4.62e-19
C701 S3 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 0.045f
C702 adder_2_0/G4 A4 0.0821f
C703 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# SUB -2.36e-19
C704 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_3_0/P3 0.00276f
C705 B3 adder_3_0/P2 8.59e-19
C706 adder_3_0/P1 A4 8.78e-20
C707 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# S4 0.0084f
C708 adder_3_0/G1 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# 0.0118f
C709 S2 CO 0.0426f
C710 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_3_0/P4 1.5e-19
C711 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# S1 3.99e-19
C712 S2 VDD 0.00253f
C713 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# CI 4.64e-20
C714 A3 A4 0.00106f
C715 adder_3_0/P1 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_47# 0.00105f
C716 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 0.00285f
C717 CO adder_2_0/sky130_fd_sc_hd__and4_1_0/a_109_47# 3.18e-19
C718 A1 adder_3_0/G2 0.00324f
C719 B3 A4 1.7f
C720 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# SUB 9.7e-20
C721 VDD adder_1_0/sky130_fd_sc_hd__and2_1_0/a_145_75# 8.07e-19
C722 SUB adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 0.00142f
C723 B4 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 0.0208f
C724 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# adder_3_0/P3 0.0039f
C725 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X adder_3_0/P3 0.00384f
C726 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# 6.41e-20
C727 adder_3_0/G1 VDD 0.694f
C728 CO adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 4.8e-20
C729 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# adder_2_0/sky130_fd_sc_hd__a21o_1_2/X -1.77e-19
C730 adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# adder_3_0/P3 0.00388f
C731 S1 adder_3_0/G3 6.53e-19
C732 VDD adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 3.32e-19
C733 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_197_47# adder_3_0/P3 4.99e-19
C734 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# CI 0.0104f
C735 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_3_0/G2 0.00133f
C736 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# B2 6.12e-20
C737 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_3_0/sky130_fd_sc_hd__xor2_1_2/B -0.014f
C738 VDD A2 0.227f
C739 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_117_297# adder_3_0/P4 9.54e-19
C740 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# adder_3_0/G1 4.07e-19
C741 adder_3_0/P3 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 1.36e-19
C742 S1 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# -1.39e-20
C743 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X adder_3_0/G3 0.0407f
C744 adder_2_0/sky130_fd_sc_hd__and4_1_0/X adder_3_0/P2 -2.14e-20
C745 B4 CI 1.51f
C746 SUB adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 9.8e-19
C747 adder_2_0/G4 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 0.0203f
C748 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# VDD 0.00935f
C749 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# A2 5.47e-19
C750 adder_3_0/G1 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# 0.00311f
C751 adder_3_0/P4 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# 2.55e-19
C752 S2 adder_3_0/P3 0.238f
C753 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X adder_3_0/G2 0.0356f
C754 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_3_0/P2 -9.82e-21
C755 adder_3_0/P1 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 0.0274f
C756 adder_2_0/G4 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 3.23e-20
C757 VDD adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# -6.01e-19
C758 S3 adder_3_0/P4 0.0135f
C759 B4 adder_3_0/P4 0.0321f
C760 adder_3_0/P3 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_109_47# 4.98e-19
C761 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# CI 2.49e-19
C762 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_117_297# adder_3_0/P4 1.04e-19
C763 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# CO 2.53e-19
C764 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 0.00297f
C765 A3 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 5.54e-20
C766 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 2.13e-20
C767 SUB CI 1.48f
C768 adder_3_0/G1 adder_3_0/P3 8.5e-20
C769 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# adder_3_0/P2 -8.74e-21
C770 B3 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 1.6e-20
C771 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# A4 0.00128f
C772 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# SUB 1.04e-19
C773 B4 B2 4.83e-19
C774 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# adder_3_0/G2 0.0051f
C775 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_3_0/P2 -1.88e-20
C776 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_3_0/P3 7.39e-20
C777 adder_2_0/G4 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_47# 6.97e-19
C778 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_3_0/P2 0.00628f
C779 A2 adder_3_0/P3 2.27e-19
C780 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# 7.13e-21
C781 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 8.3e-19
C782 SUB adder_3_0/P4 0.492f
C783 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_117_297# adder_3_0/P4 0.00227f
C784 S3 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.0023f
C785 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_384_47# adder_3_0/G2 4.16e-19
C786 CO adder_3_0/G3 4.09e-20
C787 S2 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 0.0038f
C788 adder_3_0/P1 B1 0.0278f
C789 adder_2_0/G4 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 1.75e-19
C790 VDD adder_3_0/G3 0.253f
C791 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 0 0.00137f
C792 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 0 0.255f
C793 A2 0 0.553f
C794 B2 0 0.632f
C795 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 0 0.00137f
C796 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 0 0.255f
C797 A1 0 0.469f
C798 B1 0 0.496f
C799 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0 0.00137f
C800 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 0 0.255f
C801 B4 0 1.05f
C802 A4 0 0.714f
C803 adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 0 0.177f
C804 B3 0 0.683f
C805 A3 0 0.729f
C806 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 0 0.177f
C807 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 0 0.177f
C808 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# 0 0.177f
C809 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 0 0.00137f
C810 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 0 0.255f
C811 S3 0 0.233f
C812 adder_3_0/P3 0 1.49f
C813 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 0 0.00137f
C814 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 0 0.255f
C815 SUB 0 9.62f
C816 S2 0 0.212f
C817 adder_3_0/P2 0 1.26f
C818 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 0 0.486f
C819 VDD 0 17.4f
C820 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 0 0.00137f
C821 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 0 0.255f
C822 S1 0 0.353f
C823 adder_3_0/P1 0 1.11f
C824 CI 0 2.13f
C825 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0 0.00137f
C826 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 0 0.255f
C827 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 0 0.336f
C828 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0 1.53f
C829 adder_3_0/G3 0 0.718f
C830 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 0 0.0348f
C831 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0 0.147f
C832 adder_3_0/G2 0 0.642f
C833 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 0 0.0348f
C834 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 0 0.147f
C835 adder_3_0/G1 0 0.527f
C836 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# 0 0.0348f
C837 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 0 0.147f
C838 S4 0 0.344f
C839 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 0 0.00137f
C840 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 0 0.255f
C841 adder_2_0/sky130_fd_sc_hd__and4_1_0/X 0 0.154f
C842 adder_3_0/P4 0 1.62f
C843 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 0 0.175f
C844 CO 0 0.959f
C845 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# 0 0.0348f
C846 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# 0 0.147f
C847 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 0 0.168f
C848 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 0 0.129f
C849 adder_2_0/G4 0 0.596f
C850 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 0 0.0348f
C851 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0 0.147f
C852 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 0 0.223f
C853 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 0 0.0348f
C854 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 0 0.147f
C855 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# 0 0.0348f
C856 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 0 0.147f
.ends

.subckt adder A1 B1 A2 B2 A3 B3 A4 B4 A5 B5 A6 B6 A7 B7 A8 B8 A9 B9 A10 B10 A11 B11
+ A12 B12 A13 B13 A14 B14 A15 B15 A16 B16 S1 S2 S3 S4 S5 S6 S7 S8 S9 S10 S11 S12 S13
+ S14 S15 S16 CI CO
Xadder_4_1 A5 B5 A6 B6 S5 S6 S7 S8 adder_4_2/CI adder_4_1/VDD adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75#
+ adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_384_47# adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297#
+ adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# adder_4_1/adder_2_0/sky130_fd_sc_hd__a21o_1_2/X
+ adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21#
+ adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75#
+ adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_47#
+ adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75#
+ adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297#
+ adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297#
+ adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_384_47#
+ adder_4_1/adder_2_0/sky130_fd_sc_hd__and4_1_0/X adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297#
+ adder_4_1/adder_3_0/G3 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297#
+ adder_4_1/adder_3_0/G2 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_4_1/adder_3_0/G1
+ adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297#
+ adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B
+ adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# adder_4_1/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21#
+ A8 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297#
+ adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_47# A7 adder_4_1/adder_3_0/P4
+ B8 B7 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_145_75# adder_4_1/adder_3_0/P3
+ adder_4_1/adder_3_0/P2 adder_4_1/CI adder_4_1/adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47#
+ adder_4_1/adder_3_0/P1 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297#
+ SUB adder_4_1/adder_2_0/G4 adder_4
Xadder_4_2 A9 B9 A10 B10 S9 S10 S11 S12 adder_4_3/CI adder_4_2/VDD adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75#
+ adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_384_47# adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297#
+ adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# adder_4_2/adder_2_0/sky130_fd_sc_hd__a21o_1_2/X
+ adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21#
+ adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75#
+ adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_47#
+ adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75#
+ adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297#
+ adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297#
+ adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_384_47#
+ adder_4_2/adder_2_0/sky130_fd_sc_hd__and4_1_0/X adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297#
+ adder_4_2/adder_3_0/G3 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297#
+ adder_4_2/adder_3_0/G2 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_4_2/adder_3_0/G1
+ adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297#
+ adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B
+ adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# adder_4_2/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21#
+ A12 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297#
+ adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_47# A11 adder_4_2/adder_3_0/P4
+ B12 B11 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_145_75# adder_4_2/adder_3_0/P3
+ adder_4_2/adder_3_0/P2 adder_4_2/CI adder_4_2/adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47#
+ adder_4_2/adder_3_0/P1 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297#
+ SUB adder_4_2/adder_2_0/G4 adder_4
Xadder_4_3 A13 B13 A14 B14 S13 S14 S15 S16 CO adder_4_3/VDD adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75#
+ adder_4_3/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_384_47# adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297#
+ adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# adder_4_3/adder_2_0/sky130_fd_sc_hd__a21o_1_2/X
+ adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_4_3/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21#
+ adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75#
+ adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_47#
+ adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75#
+ adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297#
+ adder_4_3/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297#
+ adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_4_3/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_384_47#
+ adder_4_3/adder_2_0/sky130_fd_sc_hd__and4_1_0/X adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297#
+ adder_4_3/adder_3_0/G3 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297#
+ adder_4_3/adder_3_0/G2 adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_4_3/adder_3_0/G1
+ adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297#
+ adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B
+ adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# adder_4_3/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21#
+ A16 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297#
+ adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_47# A15 adder_4_3/adder_3_0/P4
+ B16 B15 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_145_75# adder_4_3/adder_3_0/P3
+ adder_4_3/adder_3_0/P2 adder_4_3/CI adder_4_3/adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47#
+ adder_4_3/adder_3_0/P1 adder_4_3/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297#
+ SUB adder_4_3/adder_2_0/G4 adder_4
Xadder_4_0 A1 B1 A2 B2 S1 S2 S3 S4 adder_4_1/CI adder_4_0/VDD adder_4_0/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75#
+ adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_384_47# adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297#
+ adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# adder_4_0/adder_2_0/sky130_fd_sc_hd__a21o_1_2/X
+ adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21#
+ adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# adder_4_0/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75#
+ adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_47#
+ adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_4_0/adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75#
+ adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297#
+ adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297#
+ adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_384_47#
+ adder_4_0/adder_2_0/sky130_fd_sc_hd__and4_1_0/X adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297#
+ adder_4_0/adder_3_0/G3 adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297#
+ adder_4_0/adder_3_0/G2 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_4_0/adder_3_0/G1
+ adder_4_0/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297#
+ adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B
+ adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# adder_4_0/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21#
+ A4 adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297#
+ adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_47# A3 adder_4_0/adder_3_0/P4
+ B4 B3 adder_4_0/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_145_75# adder_4_0/adder_3_0/P3
+ adder_4_0/adder_3_0/P2 CI adder_4_0/adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47#
+ adder_4_0/adder_3_0/P1 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297#
+ SUB adder_4_0/adder_2_0/G4 adder_4
C0 adder_4_1/VDD B6 -1.33e-33
C1 B6 adder_4_1/CI 5.55e-35
C2 B7 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 2.72e-21
C3 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 3.22e-19
C4 S11 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 5.56e-20
C5 SUB adder_4_1/adder_3_0/P3 1.01e-20
C6 S3 B8 4.77e-19
C7 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_384_47# adder_4_1/adder_3_0/G1 8.69e-22
C8 A15 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 2.46e-19
C9 B16 adder_4_2/adder_3_0/P4 1.24e-19
C10 adder_4_2/adder_3_0/P4 S5 1.83e-20
C11 A14 adder_4_2/adder_3_0/G3 8.92e-19
C12 adder_4_1/adder_3_0/G2 A12 1.02e-19
C13 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_4_0/adder_3_0/P2 3.6e-19
C14 A5 CI 3.01e-20
C15 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_4_3/adder_3_0/G2 0.00265f
C16 B10 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 2.01e-20
C17 B14 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 4.05e-19
C18 B11 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 2.72e-21
C19 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# 7.69e-21
C20 adder_4_0/adder_3_0/G1 adder_4_1/CI 1.58e-19
C21 adder_4_0/adder_3_0/G1 adder_4_1/VDD 5.65e-20
C22 S3 A8 0.00571f
C23 adder_4_3/VDD adder_4_2/adder_3_0/P1 0.00122f
C24 B7 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 2.7e-20
C25 adder_4_2/CI adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 2.04e-20
C26 adder_4_1/adder_3_0/G3 adder_4_0/adder_3_0/P3 2.38e-20
C27 adder_4_2/adder_2_0/sky130_fd_sc_hd__and4_1_0/X adder_4_3/CI 3.77e-21
C28 adder_4_2/adder_3_0/G1 adder_4_1/adder_3_0/P1 7.91e-22
C29 A7 CI 2.75e-19
C30 adder_4_3/VDD adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 5.65e-20
C31 adder_4_1/adder_3_0/P1 A11 1.89e-19
C32 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 7.91e-21
C33 B8 adder_4_0/adder_3_0/G3 1.27e-19
C34 B16 A15 1.11e-34
C35 B7 adder_4_0/adder_3_0/P2 3.03e-19
C36 S3 adder_4_1/CI 7.11e-33
C37 adder_4_1/VDD S3 2.72e-19
C38 SUB adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# 1.39e-20
C39 S7 A12 0.00571f
C40 adder_4_2/VDD adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 1.01e-19
C41 A8 adder_4_0/adder_3_0/G3 1.06e-19
C42 SUB B5 1.84e-19
C43 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# A12 3.19e-20
C44 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# adder_4_0/adder_3_0/P1 2.06e-19
C45 A14 adder_4_2/adder_3_0/P1 1.27e-19
C46 A16 adder_4_2/adder_3_0/P3 4.13e-19
C47 A11 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 6.15e-20
C48 A14 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 3.9e-19
C49 B14 adder_4_2/adder_3_0/G1 7.06e-20
C50 adder_4_1/adder_3_0/G3 A11 7.8e-20
C51 adder_4_3/adder_2_0/G4 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 3.82e-21
C52 adder_4_1/VDD adder_4_0/adder_3_0/G3 5.85e-20
C53 adder_4_1/CI adder_4_0/adder_3_0/G3 1.54e-19
C54 adder_4_1/adder_3_0/P3 adder_4_2/CI 7.78e-19
C55 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_4_1/adder_3_0/G2 0.00265f
C56 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# adder_4_3/CI 3.96e-19
C57 B15 adder_4_2/adder_3_0/G3 9.04e-20
C58 A15 adder_4_2/adder_3_0/P3 2.29e-19
C59 A16 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 4.77e-20
C60 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# S8 2.71e-19
C61 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# S9 5.99e-21
C62 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_4_0/adder_3_0/P3 1.33e-20
C63 adder_4_0/adder_3_0/G2 A7 7.47e-20
C64 S10 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 2.19e-20
C65 A15 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 3.5e-20
C66 A16 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 1.39e-19
C67 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 7.69e-21
C68 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B A13 1.22e-19
C69 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# adder_4_2/CI 9.5e-20
C70 adder_4_2/adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# adder_4_3/CI 2.13e-21
C71 SUB adder_4_2/CI 0.04f
C72 B12 adder_4_1/adder_3_0/G1 1.31e-19
C73 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# S5 5.99e-21
C74 A15 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 6.15e-20
C75 adder_4_2/adder_3_0/P1 B15 2.28e-19
C76 B16 S10 3.18e-19
C77 SUB A6 4.78e-19
C78 S1 B8 2.42e-19
C79 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# B15 2.7e-20
C80 S11 adder_4_3/CI 7.11e-33
C81 adder_4_0/adder_3_0/P4 B8 1.24e-19
C82 S1 A8 1.3e-19
C83 A16 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 3.39e-20
C84 B12 adder_4_1/adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 1.9e-21
C85 S1 adder_4_1/CI 2.87e-19
C86 S1 adder_4_1/VDD 8.75e-19
C87 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# A10 1.76e-20
C88 adder_4_0/adder_3_0/P4 adder_4_1/VDD 1.01e-19
C89 A10 adder_4_1/VDD 2.23e-20
C90 A10 adder_4_1/CI 1.92e-19
C91 B12 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 3.74e-19
C92 adder_4_2/adder_3_0/P1 B13 8.38e-20
C93 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# A7 2.46e-19
C94 SUB S12 6.99e-20
C95 S4 B8 5.46e-19
C96 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# B10 2.01e-20
C97 A11 adder_4_1/adder_3_0/G1 8.1e-20
C98 adder_4_2/adder_3_0/G2 adder_4_3/CI 1.47e-19
C99 adder_4_3/VDD adder_4_3/CI 0.0264f
C100 B10 adder_4_1/VDD 2.46e-19
C101 B10 adder_4_1/CI 8.69e-19
C102 B14 A13 1.11e-34
C103 A16 adder_4_2/adder_3_0/P2 3.39e-19
C104 A8 S4 3.33e-19
C105 adder_4_1/adder_3_0/P3 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 1.33e-20
C106 adder_4_1/adder_3_0/P3 adder_4_2/adder_3_0/P3 1.88e-19
C107 adder_4_1/adder_3_0/G2 CI 8.7e-21
C108 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# A7 3.5e-20
C109 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 3.19e-22
C110 SUB B16 0.00215f
C111 adder_4_1/adder_3_0/P2 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 5.27e-22
C112 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 6.83e-22
C113 B9 adder_4_1/adder_3_0/G2 1.61e-19
C114 adder_4_3/VDD S11 2.72e-19
C115 S9 adder_4_3/CI 2.87e-19
C116 B7 adder_4_0/VDD 4.79e-20
C117 A15 adder_4_2/adder_3_0/P2 1.97e-19
C118 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B B5 4.08e-21
C119 adder_4_1/VDD S4 2.91e-19
C120 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_1/adder_3_0/P2 2.19e-20
C121 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# A12 3.19e-20
C122 B10 B11 4.44e-34
C123 B6 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 2.01e-20
C124 B6 adder_4_0/adder_3_0/P3 0.00256f
C125 adder_4_1/VDD A12 6.31e-20
C126 adder_4_1/CI A12 5.12e-19
C127 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# adder_4_2/VDD 4.75e-20
C128 SUB adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 1.39e-20
C129 adder_4_3/VDD adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 5.51e-20
C130 adder_4_3/adder_3_0/G1 adder_4_2/adder_3_0/P1 7.91e-22
C131 adder_4_2/adder_3_0/P1 adder_4_1/CI 2.44e-20
C132 A10 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 2.29e-19
C133 SUB adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 1.66e-20
C134 A11 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 2.34e-20
C135 SUB adder_4_2/adder_3_0/P3 1.01e-20
C136 B7 adder_4_0/adder_3_0/G1 9.39e-20
C137 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B B8 0.00191f
C138 B10 adder_4_2/VDD 5.55e-32
C139 adder_4_2/adder_3_0/G3 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 3.18e-20
C140 B10 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 4.05e-19
C141 SUB adder_4_1/adder_2_0/G4 4.83e-20
C142 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B A8 0.0011f
C143 adder_4_3/adder_2_0/G4 adder_4_3/CI 3.53e-20
C144 adder_4_3/VDD adder_4_2/adder_3_0/G2 3.95e-20
C145 S1 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 6.6e-21
C146 adder_4_3/adder_3_0/P3 S10 1.88e-20
C147 B16 adder_4_2/CI 7.74e-19
C148 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_1/adder_3_0/P1 4.66e-20
C149 adder_4_2/CI S5 2.87e-19
C150 A7 B8 1.11e-34
C151 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 5.8e-21
C152 SUB adder_4_3/adder_3_0/G3 5.02e-20
C153 B15 adder_4_3/CI 7.76e-19
C154 S11 adder_4_3/adder_2_0/G4 2.25e-20
C155 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_4_1/CI 0.433f
C156 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_4_1/VDD 0.00127f
C157 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_4_3/CI 2.04e-20
C158 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 7.91e-21
C159 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_4_0/adder_3_0/G3 2.84e-32
C160 adder_4_3/VDD S9 8.75e-19
C161 A14 adder_4_2/adder_3_0/G2 5.72e-20
C162 SUB adder_4_1/adder_3_0/P2 4.74e-20
C163 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B A6 4.4e-20
C164 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_4_2/CI 1.52e-20
C165 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B A12 0.0011f
C166 S8 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 7.81e-20
C167 A7 adder_4_1/CI 0.00338f
C168 B7 adder_4_0/adder_3_0/G3 9.04e-20
C169 A16 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 3.19e-20
C170 adder_4_2/adder_3_0/P1 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 2.81e-20
C171 adder_4_2/adder_2_0/G4 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 9.08e-21
C172 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# A13 2.68e-19
C173 adder_4_2/CI adder_4_2/adder_3_0/P3 3.24e-20
C174 adder_4_2/CI adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 2.86e-20
C175 adder_4_1/CI adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 2.04e-20
C176 S8 adder_4_2/VDD 2.91e-19
C177 S12 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 7.81e-20
C178 B5 adder_4_0/adder_3_0/P1 8.38e-20
C179 SUB adder_4_0/adder_3_0/P1 -1.14e-31
C180 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 3.52e-21
C181 A15 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 2.32e-20
C182 B16 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 5.68e-20
C183 adder_4_2/CI adder_4_1/adder_2_0/G4 1.64e-21
C184 B15 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 2.9e-20
C185 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# A6 1.76e-20
C186 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 3.2e-20
C187 B16 S12 5.46e-19
C188 adder_4_1/adder_3_0/P3 adder_4_2/adder_3_0/P2 2.36e-20
C189 S6 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 5.48e-20
C190 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 7.91e-21
C191 SUB adder_4_3/adder_3_0/P3 1.01e-20
C192 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_4_3/CI 4.64e-20
C193 adder_4_1/CI adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 2.8e-20
C194 B12 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 2.14e-19
C195 B5 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 1.56e-20
C196 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 6.83e-22
C197 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 3.2e-20
C198 adder_4_2/CI adder_4_1/adder_3_0/P2 9.44e-19
C199 B15 adder_4_2/adder_3_0/G2 8.67e-20
C200 adder_4_3/VDD B15 5.68e-32
C201 adder_4_3/adder_2_0/G4 S9 1.75e-20
C202 SUB adder_4_0/adder_3_0/P2 -5.68e-32
C203 SUB adder_4_1/adder_3_0/G3 5.02e-20
C204 SUB adder_4_3/adder_3_0/G2 1.6e-20
C205 SUB B14 6.79e-19
C206 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# A9 2.25e-19
C207 B8 CI 7.74e-19
C208 SUB adder_4_2/adder_3_0/P2 4.74e-20
C209 adder_4_1/VDD A9 7.39e-21
C210 adder_4_1/CI A9 3.01e-20
C211 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# B11 4.06e-20
C212 S9 B15 8.93e-20
C213 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 3.52e-21
C214 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# S9 5.99e-21
C215 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 1.42e-19
C216 A8 CI 5.12e-19
C217 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# S5 5.99e-21
C218 A6 adder_4_0/adder_3_0/P1 1.27e-19
C219 B16 adder_4_2/adder_3_0/P3 5.72e-19
C220 adder_4_2/adder_3_0/P3 S5 1.67e-20
C221 B7 S1 8.93e-20
C222 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# adder_4_1/adder_2_0/G4 3.82e-21
C223 adder_4_2/CI adder_4_1/adder_3_0/P1 4.71e-19
C224 A6 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 1.53e-19
C225 adder_4_1/adder_3_0/P4 adder_4_1/CI 3.66e-20
C226 S2 A7 3.71e-20
C227 S2 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 1.18e-20
C228 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_4_2/VDD 5.65e-20
C229 adder_4_1/CI CI 0.0496f
C230 adder_4_1/VDD CI 9.52e-19
C231 B13 adder_4_2/adder_3_0/G2 1.61e-19
C232 B16 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 5.68e-20
C233 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# B11 4.21e-20
C234 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# B9 1.56e-20
C235 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 9.13e-20
C236 adder_4_2/adder_3_0/P1 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 2.06e-19
C237 B9 adder_4_1/VDD 5.18e-20
C238 B9 adder_4_1/CI 1.09e-19
C239 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_4_3/VDD 5.65e-20
C240 adder_4_2/CI adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 2.02e-19
C241 SUB adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 1.66e-20
C242 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# A6 1.76e-20
C243 adder_4_2/CI adder_4_1/adder_3_0/G3 1.54e-19
C244 B16 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 1.66e-19
C245 adder_4_2/CI adder_4_3/adder_3_0/G2 8.7e-21
C246 adder_4_2/adder_3_0/P3 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 3.3e-19
C247 B12 S8 5.46e-19
C248 B14 adder_4_2/CI 8.69e-19
C249 SUB adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 1.39e-20
C250 adder_4_0/adder_3_0/G2 B8 1.21e-19
C251 A6 adder_4_0/adder_3_0/P2 1.62e-19
C252 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_2/VDD 4.95e-20
C253 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B A9 3.79e-20
C254 adder_4_0/adder_3_0/G2 A8 1.02e-19
C255 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# A14 1.76e-20
C256 adder_4_2/VDD adder_4_3/CI 0.00644f
C257 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 6.83e-22
C258 adder_4_2/VDD adder_4_1/adder_3_0/P4 1.01e-19
C259 B11 S6 3.58e-19
C260 adder_4_1/adder_3_0/G2 adder_4_1/CI 6.94e-36
C261 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 6.83e-22
C262 adder_4_2/adder_3_0/G2 adder_4_1/CI 8.7e-21
C263 adder_4_0/adder_3_0/G2 adder_4_1/CI 1.47e-19
C264 adder_4_0/adder_3_0/G2 adder_4_1/VDD 3.95e-20
C265 adder_4_3/adder_3_0/G1 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_384_47# 8.69e-22
C266 adder_4_3/VDD adder_4_3/adder_3_0/G1 2.84e-32
C267 adder_4_2/adder_3_0/P3 adder_4_3/adder_3_0/G3 2.38e-20
C268 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# B11 2.9e-20
C269 S7 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_145_75# 1.39e-20
C270 adder_4_3/CI adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 5.9e-20
C271 adder_4_2/adder_3_0/G1 A12 -1.39e-35
C272 S6 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 2.19e-20
C273 adder_4_2/adder_2_0/G4 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 3.82e-21
C274 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# CI 5.01e-20
C275 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_4_1/adder_3_0/P2 2.53e-19
C276 SUB adder_4_1/adder_3_0/G1 6.38e-21
C277 B9 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.00399f
C278 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 9.13e-20
C279 SUB adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 1.39e-20
C280 adder_4_2/VDD S6 3.45e-19
C281 B8 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 5.68e-20
C282 B11 adder_4_1/adder_3_0/G2 8.67e-20
C283 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_4_2/VDD 5.51e-20
C284 S2 adder_4_1/adder_3_0/P4 2.06e-20
C285 B11 adder_4_2/adder_3_0/G2 1.39e-35
C286 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# S4 2.71e-19
C287 A8 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 3.71e-19
C288 adder_4_3/adder_3_0/G3 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 6.86e-21
C289 B7 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.00977f
C290 B8 adder_4_0/adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 1.9e-21
C291 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# B15 2.7e-20
C292 A7 adder_4_0/adder_3_0/P3 2.29e-19
C293 A7 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 2.32e-20
C294 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# B8 5.68e-20
C295 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# S10 1.82e-19
C296 S2 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# 1.82e-19
C297 B16 adder_4_2/adder_3_0/P2 4.43e-19
C298 adder_4_2/VDD adder_4_1/adder_3_0/G2 3.95e-20
C299 adder_4_1/VDD adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 5.51e-20
C300 adder_4_3/adder_3_0/P4 adder_4_3/CI 3.66e-20
C301 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# A8 4.77e-20
C302 B12 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 5.68e-20
C303 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_4_1/adder_3_0/G3 6.86e-21
C304 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_4_1/adder_2_0/G4 9.08e-21
C305 adder_4_2/adder_3_0/P3 adder_4_3/adder_3_0/P3 1.88e-19
C306 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# B11 2.7e-20
C307 adder_4_2/adder_3_0/G2 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.00265f
C308 B5 adder_4_0/VDD 5.18e-20
C309 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# B8 5.68e-20
C310 S7 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 2.47e-20
C311 adder_4_2/CI adder_4_1/adder_3_0/G1 1.58e-19
C312 S11 adder_4_3/adder_3_0/P4 2.35e-20
C313 adder_4_1/CI adder_4_0/adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 2.13e-21
C314 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 4.28e-21
C315 adder_4_3/VDD adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 1.01e-19
C316 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# A8 4.77e-20
C317 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_1/CI 7.44e-19
C318 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_1/VDD 4.95e-20
C319 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_4_2/adder_3_0/P2 1.18e-20
C320 SUB B6 6.79e-19
C321 adder_4_3/adder_3_0/G2 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_384_47# 4.9e-21
C322 S7 adder_4_2/VDD 2.72e-19
C323 adder_4_1/adder_3_0/P2 adder_4_0/adder_3_0/P1 1.07e-21
C324 A14 adder_4_2/VDD 2.23e-20
C325 adder_4_2/adder_3_0/P3 adder_4_3/adder_3_0/G2 3.43e-21
C326 A16 adder_4_2/adder_3_0/G3 1.06e-19
C327 B14 adder_4_2/adder_3_0/P3 0.00256f
C328 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_4_2/VDD 5.65e-20
C329 B12 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 5.68e-20
C330 B16 adder_4_2/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# 2.93e-22
C331 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# B13 1.56e-20
C332 B5 adder_4_0/adder_3_0/G1 5.49e-20
C333 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 9.13e-20
C334 A16 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 6.43e-20
C335 SUB adder_4_0/adder_3_0/G1 5.68e-32
C336 adder_4_3/adder_3_0/P2 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 3.15e-20
C337 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_4_1/VDD 5.65e-20
C338 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_4_1/CI 6.87e-20
C339 A15 adder_4_2/adder_3_0/G3 7.8e-20
C340 adder_4_2/CI adder_4_1/adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 2.13e-21
C341 B14 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 2.06e-22
C342 A14 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 1.53e-19
C343 B12 adder_4_1/adder_3_0/P4 1.24e-19
C344 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# S10 5.48e-20
C345 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 4.28e-21
C346 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_4_3/CI 0.433f
C347 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 5e-21
C348 B14 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 5.78e-20
C349 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# A11 3.5e-20
C350 A16 adder_4_2/adder_3_0/P1 2.81e-19
C351 adder_4_2/CI adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 5.9e-20
C352 adder_4_3/adder_3_0/G3 adder_4_2/adder_3_0/P2 4e-21
C353 adder_4_1/adder_3_0/P2 adder_4_0/adder_3_0/P2 2.08e-20
C354 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# S3 2.47e-20
C355 A8 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 3.39e-20
C356 adder_4_2/adder_3_0/P1 A13 2.83e-20
C357 A10 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 1.76e-20
C358 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# A12 3.39e-20
C359 adder_4_0/VDD A6 2.23e-20
C360 A16 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 3.19e-20
C361 adder_4_2/adder_3_0/P4 S8 2.69e-20
C362 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# CI 2.8e-20
C363 B12 S6 3.18e-19
C364 adder_4_2/adder_3_0/P2 adder_4_1/adder_3_0/P2 2.08e-20
C365 B12 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 5.68e-20
C366 SUB adder_4_0/adder_3_0/G3 -1.42e-32
C367 B15 adder_4_2/VDD 4.79e-20
C368 A15 adder_4_2/adder_3_0/P1 1.89e-19
C369 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# 7.69e-21
C370 adder_4_3/adder_2_0/G4 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 9.08e-21
C371 B10 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 2.01e-20
C372 S9 adder_4_3/adder_3_0/P4 1.83e-20
C373 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# adder_4_1/CI 9.5e-20
C374 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# CI 9.5e-20
C375 B16 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 3.81e-20
C376 A15 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 2.32e-20
C377 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# A11 2.46e-19
C378 B7 CI 3.65e-19
C379 adder_4_1/VDD B8 -1.11e-34
C380 B8 adder_4_1/CI 0.279f
C381 adder_4_2/adder_3_0/G1 adder_4_3/CI 1.58e-19
C382 B16 adder_4_2/adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 4.4e-21
C383 adder_4_0/adder_3_0/G1 A6 6.2e-20
C384 B15 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 2.72e-21
C385 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 5.92e-22
C386 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 3.52e-21
C387 adder_4_1/adder_3_0/P1 adder_4_0/adder_3_0/P2 0.00296f
C388 B12 adder_4_1/adder_3_0/G2 1.21e-19
C389 A8 adder_4_1/CI 0.00128f
C390 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 7.91e-21
C391 adder_4_2/adder_3_0/P2 adder_4_1/adder_3_0/P1 1.07e-21
C392 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# A12 3.19e-20
C393 SUB adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 1.17e-20
C394 adder_4_3/VDD adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.00127f
C395 adder_4_1/adder_3_0/P3 S1 1.67e-20
C396 adder_4_1/VDD adder_4_1/CI 0.0264f
C397 SUB adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 1.39e-20
C398 B13 adder_4_2/VDD 5.18e-20
C399 adder_4_1/adder_3_0/P3 A10 4.46e-20
C400 adder_4_1/adder_3_0/G3 adder_4_0/adder_3_0/P2 4e-21
C401 B12 S7 4.77e-19
C402 adder_4_1/adder_3_0/G2 adder_4_0/adder_3_0/P3 3.43e-21
C403 A11 S6 3.71e-20
C404 adder_4_1/adder_3_0/P1 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 2.06e-19
C405 B12 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 3.81e-20
C406 B7 adder_4_1/adder_3_0/G2 1.39e-35
C407 adder_4_2/adder_3_0/P2 adder_4_3/adder_3_0/G2 6.64e-21
C408 B14 adder_4_2/adder_3_0/P2 1.84e-19
C409 A6 adder_4_0/adder_3_0/G3 8.92e-19
C410 adder_4_1/adder_3_0/P3 adder_4_2/adder_3_0/G3 2.38e-20
C411 B7 adder_4_0/adder_3_0/G2 8.67e-20
C412 A14 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 2.29e-19
C413 adder_4_1/adder_3_0/P3 B10 0.00256f
C414 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 5.92e-22
C415 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# CI 2.46e-19
C416 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_4_0/adder_3_0/P1 5.99e-21
C417 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# B11 2.7e-20
C418 adder_4_1/VDD B11 4.79e-20
C419 B11 adder_4_1/CI 3.65e-19
C420 adder_4_2/adder_2_0/G4 adder_4_3/CI 1.64e-21
C421 adder_4_2/adder_2_0/G4 adder_4_1/adder_3_0/P4 3.69e-21
C422 A11 adder_4_1/adder_3_0/G2 7.47e-20
C423 adder_4_3/VDD adder_4_2/adder_3_0/G1 5.65e-20
C424 SUB A10 4.78e-19
C425 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B B6 5.78e-20
C426 adder_4_2/CI adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_47# 8.76e-20
C427 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# S1 6.6e-21
C428 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 5.92e-22
C429 adder_4_1/adder_3_0/P2 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 1.18e-20
C430 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_4_2/VDD 5.65e-20
C431 adder_4_1/adder_3_0/P3 A12 4.13e-19
C432 adder_4_2/VDD adder_4_1/CI 9.52e-19
C433 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_4_0/adder_3_0/P2 2.53e-19
C434 SUB adder_4_2/adder_3_0/G3 5.02e-20
C435 S2 B8 3.18e-19
C436 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# S10 1.18e-20
C437 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_2/CI 5.01e-20
C438 SUB B10 6.79e-19
C439 adder_4_2/adder_2_0/G4 S6 1.98e-20
C440 A14 adder_4_2/adder_3_0/G1 6.2e-20
C441 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_4_0/adder_3_0/P2 1.18e-20
C442 adder_4_0/adder_3_0/P1 adder_4_1/adder_3_0/G1 7.91e-22
C443 S2 A8 1.69e-19
C444 B7 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 2.9e-20
C445 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# B6 2.01e-20
C446 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# A11 2.32e-20
C447 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B B15 0.00977f
C448 A16 adder_4_3/CI 0.00128f
C449 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 1.75e-20
C450 B11 adder_4_2/VDD 5.68e-32
C451 SUB S4 6.99e-20
C452 adder_4_1/adder_3_0/P1 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 5.99e-21
C453 S2 adder_4_1/CI 0.0018f
C454 B11 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.00977f
C455 SUB A12 0.00154f
C456 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_4_1/CI 3.7e-20
C457 S2 adder_4_1/VDD 3.45e-19
C458 adder_4_2/CI adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 1.39e-35
C459 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# S4 7.81e-20
C460 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# B7 4.21e-20
C461 A15 adder_4_3/CI 0.00338f
C462 S11 A16 0.00571f
C463 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 7.91e-21
C464 adder_4_2/adder_3_0/P4 S6 2.06e-20
C465 adder_4_1/adder_3_0/P3 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 1.97e-20
C466 SUB S8 6.99e-20
C467 S3 adder_4_1/adder_2_0/G4 2.25e-20
C468 B14 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 2.01e-20
C469 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_47# S12 1.16e-19
C470 adder_4_2/CI B10 5.55e-35
C471 adder_4_2/CI adder_4_2/adder_3_0/G3 4.85e-20
C472 adder_4_2/VDD adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.00127f
C473 B7 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 4.06e-20
C474 A16 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 3.71e-19
C475 adder_4_2/adder_3_0/G1 B15 9.39e-20
C476 S7 adder_4_2/adder_2_0/G4 2.25e-20
C477 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# A9 2.68e-19
C478 B13 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.00399f
C479 SUB adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 1.76e-20
C480 B6 adder_4_0/adder_3_0/P1 1.48e-19
C481 B6 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 2.79e-20
C482 adder_4_3/VDD adder_4_2/adder_3_0/P4 1.01e-19
C483 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B B5 0.00399f
C484 SUB A5 1.99e-19
C485 SUB adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 3.41e-20
C486 A16 adder_4_2/adder_3_0/G2 1.02e-19
C487 adder_4_2/CI A12 0.00128f
C488 B12 adder_4_1/adder_2_0/sky130_fd_sc_hd__and4_1_0/X 3.37e-21
C489 SUB A7 8.93e-19
C490 S6 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# 1.82e-19
C491 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# B12 3.81e-20
C492 SUB adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 1.76e-20
C493 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# B6 2.01e-20
C494 A15 adder_4_2/adder_3_0/G2 7.47e-20
C495 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# B8 3.81e-20
C496 B8 adder_4_0/adder_3_0/P3 5.72e-19
C497 adder_4_2/adder_3_0/P4 S7 2.35e-20
C498 B12 adder_4_1/VDD 6.98e-19
C499 B12 adder_4_1/CI 7.74e-19
C500 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 5.8e-21
C501 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_4_2/adder_3_0/P3 3.44e-19
C502 adder_4_3/CI S10 0.0018f
C503 A16 S9 1.3e-19
C504 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_2/adder_3_0/P3 2.47e-20
C505 adder_4_2/adder_3_0/G1 B13 5.49e-20
C506 B7 B8 2.22e-34
C507 B6 adder_4_0/adder_3_0/P2 1.84e-19
C508 A8 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 3.19e-20
C509 A8 adder_4_0/adder_3_0/P3 4.13e-19
C510 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_4_3/adder_3_0/P1 2.81e-20
C511 S2 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 5.48e-20
C512 A15 S9 1.1e-19
C513 B16 adder_4_2/adder_3_0/G3 1.27e-19
C514 adder_4_2/adder_3_0/G3 S5 1.85e-20
C515 adder_4_1/CI adder_4_0/adder_3_0/P3 7.78e-19
C516 adder_4_1/VDD adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 5.65e-20
C517 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_4_1/CI 4.64e-20
C518 adder_4_1/VDD adder_4_0/adder_3_0/P3 0.00144f
C519 SUB adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 1.01e-20
C520 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# S6 1.18e-20
C521 B16 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 2.14e-19
C522 B7 adder_4_1/VDD 5.68e-32
C523 B7 adder_4_1/CI 7.44e-19
C524 adder_4_3/adder_2_0/G4 adder_4_2/adder_3_0/P4 3.69e-21
C525 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B A6 2.29e-19
C526 B12 adder_4_2/VDD -1.11e-34
C527 S1 adder_4_1/adder_2_0/G4 1.75e-20
C528 SUB adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 1.01e-20
C529 SUB adder_4_3/adder_3_0/P2 4.74e-20
C530 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# A11 2.32e-20
C531 adder_4_2/adder_3_0/G1 adder_4_1/CI 0.0031f
C532 S5 A12 1.3e-19
C533 adder_4_0/adder_3_0/P4 adder_4_1/adder_2_0/G4 3.69e-21
C534 B12 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.00191f
C535 adder_4_1/VDD A11 2.34e-19
C536 A11 adder_4_1/CI 2.75e-19
C537 SUB A9 1.99e-19
C538 B16 adder_4_2/adder_3_0/P1 3.59e-19
C539 adder_4_3/VDD S10 3.45e-19
C540 B16 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 3.81e-20
C541 SUB adder_4_3/CI 0.04f
C542 B8 adder_4_0/adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 4.4e-21
C543 SUB CI 3.79e-20
C544 B5 CI 1.09e-19
C545 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_4_2/adder_3_0/P1 5.99e-21
C546 A10 adder_4_1/adder_3_0/P2 1.62e-19
C547 adder_4_2/CI adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 6.87e-20
C548 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_0/adder_3_0/P3 2.47e-20
C549 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# 1.42e-19
C550 S7 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 5.56e-20
C551 SUB B9 1.84e-19
C552 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 7.69e-21
C553 adder_4_2/CI adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 3.96e-19
C554 adder_4_1/adder_3_0/P3 adder_4_2/adder_3_0/G2 3.43e-21
C555 B10 adder_4_1/adder_3_0/P2 1.84e-19
C556 adder_4_1/adder_3_0/P2 adder_4_2/adder_3_0/G3 4e-21
C557 SUB S6 3.33e-22
C558 adder_4_2/CI adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 2.8e-20
C559 adder_4_2/adder_3_0/G1 adder_4_2/VDD 2.84e-32
C560 adder_4_1/CI adder_4_0/adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 1.34e-20
C561 A16 B13 5.55e-35
C562 adder_4_2/CI adder_4_3/adder_3_0/P2 4.97e-20
C563 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_4_0/adder_3_0/P3 3.44e-19
C564 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B A11 4.82e-19
C565 adder_4_2/CI adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 7.44e-19
C566 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# A16 3.19e-20
C567 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# A13 2.25e-19
C568 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B A5 1.22e-19
C569 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_2/adder_3_0/P2 2.19e-20
C570 adder_4_2/adder_3_0/G1 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_384_47# 8.69e-22
C571 S2 B7 3.58e-19
C572 A10 adder_4_1/adder_3_0/P1 1.27e-19
C573 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 5e-21
C574 adder_4_0/adder_3_0/P2 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 5.27e-22
C575 adder_4_2/CI adder_4_3/CI 0.0496f
C576 adder_4_3/adder_2_0/G4 S10 1.98e-20
C577 SUB adder_4_1/adder_3_0/G2 1.6e-20
C578 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# A15 2.32e-20
C579 B16 adder_4_2/adder_2_0/sky130_fd_sc_hd__and4_1_0/X 3.37e-21
C580 adder_4_1/adder_3_0/P2 A12 3.39e-19
C581 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B A7 6.15e-20
C582 B5 adder_4_0/adder_3_0/G2 1.61e-19
C583 SUB adder_4_2/adder_3_0/G2 1.6e-20
C584 SUB adder_4_3/VDD 0.0884f
C585 adder_4_2/adder_3_0/P1 adder_4_1/adder_3_0/P2 0.00296f
C586 B10 adder_4_1/adder_3_0/P1 1.48e-19
C587 S1 adder_4_1/adder_3_0/G3 1.85e-20
C588 A10 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 4.4e-20
C589 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# A5 2.68e-19
C590 A6 CI 1.92e-19
C591 B15 S10 3.58e-19
C592 A10 adder_4_1/adder_3_0/G3 8.92e-19
C593 adder_4_0/VDD B6 2.46e-19
C594 adder_4_2/CI S6 0.0018f
C595 adder_4_3/adder_3_0/G1 A16 -1.39e-35
C596 adder_4_2/adder_3_0/G3 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 6.86e-21
C597 SUB A14 4.78e-19
C598 B10 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 5.78e-20
C599 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# A7 2.32e-20
C600 B10 adder_4_1/adder_3_0/G3 6.79e-20
C601 B14 adder_4_2/adder_3_0/G3 6.79e-20
C602 adder_4_1/adder_3_0/P1 A12 2.81e-19
C603 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_3/CI 7.44e-19
C604 adder_4_3/CI adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 3.7e-20
C605 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_4_1/adder_3_0/P2 3.15e-20
C606 adder_4_0/adder_3_0/G1 B6 7.06e-20
C607 adder_4_2/CI adder_4_1/adder_3_0/G2 1.47e-19
C608 adder_4_2/CI adder_4_2/adder_3_0/G2 6.94e-36
C609 adder_4_3/VDD adder_4_2/CI 9.52e-19
C610 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B A12 1.39e-19
C611 S1 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 5.99e-21
C612 adder_4_1/adder_3_0/P3 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 3.44e-19
C613 adder_4_1/adder_3_0/G3 A12 1.06e-19
C614 S11 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 2.47e-20
C615 adder_4_0/adder_3_0/G2 A6 5.72e-20
C616 B16 adder_4_3/CI 0.279f
C617 SUB adder_4_3/adder_2_0/G4 4.83e-20
C618 B16 adder_4_2/adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 1.9e-21
C619 A5 adder_4_0/adder_3_0/P1 2.83e-20
C620 adder_4_2/adder_3_0/P1 adder_4_3/adder_3_0/G2 5.87e-21
C621 B14 adder_4_2/adder_3_0/P1 1.48e-19
C622 A16 adder_4_2/VDD 6.31e-20
C623 A13 adder_4_2/VDD 7.39e-21
C624 B12 adder_4_2/adder_3_0/G1 -6.94e-36
C625 B14 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 2.01e-20
C626 adder_4_2/CI S7 7.11e-33
C627 A14 adder_4_2/CI 1.92e-19
C628 SUB B15 0.00112f
C629 B16 S11 4.77e-19
C630 B12 A11 1.11e-34
C631 adder_4_3/adder_3_0/P2 adder_4_2/adder_3_0/P3 2.36e-20
C632 A7 adder_4_0/adder_3_0/P1 1.89e-19
C633 SUB adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 1.66e-20
C634 adder_4_2/CI adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 4.64e-20
C635 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_4_1/adder_3_0/P1 2.81e-20
C636 B7 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 2.7e-20
C637 B7 adder_4_0/adder_3_0/P3 2.06e-19
C638 A15 adder_4_2/VDD 2.34e-19
C639 A7 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 2.34e-20
C640 A16 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 1.4e-20
C641 B6 adder_4_0/adder_3_0/G3 6.79e-20
C642 SUB adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 1.17e-20
C643 adder_4_1/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# B12 2.93e-22
C644 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 6.83e-22
C645 adder_4_2/adder_3_0/P3 adder_4_3/CI 7.78e-19
C646 A5 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 2.25e-19
C647 B16 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 5.68e-20
C648 adder_4_1/adder_3_0/P2 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 3.6e-19
C649 adder_4_3/VDD adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 4.95e-20
C650 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# B11 2.7e-20
C651 A15 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 2.34e-20
C652 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_4_1/adder_3_0/G3 3.18e-20
C653 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# A7 2.32e-20
C654 adder_4_3/VDD S12 2.91e-19
C655 A10 adder_4_1/adder_3_0/G1 6.2e-20
C656 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_4_3/CI 6.87e-20
C657 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_1/CI 5.01e-20
C658 A7 adder_4_0/adder_3_0/P2 1.97e-19
C659 B16 adder_4_2/adder_3_0/G2 1.21e-19
C660 SUB B13 1.84e-19
C661 B16 adder_4_3/VDD -1.11e-34
C662 adder_4_2/adder_3_0/P3 S6 1.88e-20
C663 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_4_2/VDD 2.78e-20
C664 B10 adder_4_1/adder_3_0/G1 7.06e-20
C665 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# 7.69e-21
C666 adder_4_3/adder_3_0/G3 adder_4_3/CI 4.85e-20
C667 S9 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 6.6e-21
C668 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_4_3/CI 2.56e-19
C669 adder_4_2/CI B15 3.65e-19
C670 SUB adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# 1.39e-20
C671 adder_4_1/adder_3_0/P1 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 6.6e-21
C672 adder_4_1/adder_3_0/P3 adder_4_1/CI 3.24e-20
C673 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_384_47# adder_4_2/adder_3_0/G2 4.9e-21
C674 SUB B8 0.00215f
C675 adder_4_2/CI adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 3.7e-20
C676 B16 S9 2.42e-19
C677 adder_4_1/adder_3_0/P2 CI 4.97e-20
C678 B5 A8 5.55e-35
C679 SUB A8 0.00154f
C680 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# adder_4_0/adder_3_0/P3 3.3e-19
C681 adder_4_1/adder_3_0/G1 A12 1.1e-19
C682 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 1.75e-20
C683 A10 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 1.53e-19
C684 adder_4_3/VDD adder_4_2/adder_3_0/P3 0.00144f
C685 adder_4_1/adder_3_0/P1 A9 2.83e-20
C686 B12 adder_4_1/adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 4.4e-21
C687 adder_4_1/adder_3_0/P3 B11 2.06e-19
C688 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 3.22e-19
C689 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 3.2e-20
C690 SUB adder_4_1/CI 0.04f
C691 SUB adder_4_1/VDD 0.0884f
C692 SUB adder_4_3/adder_3_0/G1 6.38e-21
C693 B10 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 2.79e-20
C694 adder_4_3/VDD adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 5.65e-20
C695 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_47# S8 1.16e-19
C696 adder_4_2/CI B13 1.09e-19
C697 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# B15 4.21e-20
C698 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_47# S4 1.16e-19
C699 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# adder_4_1/CI 3.7e-20
C700 adder_4_3/adder_3_0/P3 adder_4_3/CI 3.24e-20
C701 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B A9 1.22e-19
C702 A14 adder_4_2/adder_3_0/P3 4.46e-20
C703 adder_4_1/adder_3_0/P3 adder_4_2/VDD 0.00144f
C704 adder_4_1/adder_3_0/P1 CI 2.44e-20
C705 A16 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.0011f
C706 adder_4_2/adder_3_0/P2 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 3.6e-19
C707 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B A13 3.79e-20
C708 adder_4_3/adder_3_0/P2 adder_4_2/adder_3_0/P2 2.08e-20
C709 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# adder_4_1/CI 3.96e-19
C710 adder_4_3/VDD adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 1.51e-19
C711 B9 adder_4_1/adder_3_0/P1 8.38e-20
C712 SUB B11 0.00112f
C713 adder_4_1/adder_3_0/P2 adder_4_2/adder_3_0/G2 6.64e-21
C714 adder_4_3/adder_3_0/G2 adder_4_3/CI 6.94e-36
C715 B14 adder_4_3/CI 5.55e-35
C716 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B A12 1.4e-20
C717 A15 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 4.82e-19
C718 adder_4_2/adder_3_0/P2 adder_4_3/CI 6.08e-19
C719 adder_4_3/adder_3_0/G3 S9 1.85e-20
C720 adder_4_2/CI adder_4_1/adder_2_0/sky130_fd_sc_hd__and4_1_0/X 3.77e-21
C721 B9 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 4.08e-21
C722 S5 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 6.6e-21
C723 adder_4_3/adder_3_0/P4 S10 2.06e-20
C724 A14 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 4.4e-20
C725 adder_4_1/adder_3_0/G2 adder_4_0/adder_3_0/P1 5.87e-21
C726 S2 adder_4_1/adder_3_0/P3 1.88e-20
C727 adder_4_2/CI adder_4_3/adder_3_0/P1 2.44e-20
C728 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_4_2/CI 4.64e-20
C729 SUB adder_4_2/VDD 0.0884f
C730 adder_4_3/adder_3_0/G1 adder_4_2/CI 0.0031f
C731 adder_4_2/CI adder_4_1/VDD 0.00644f
C732 adder_4_2/CI adder_4_1/CI 0.0496f
C733 SUB adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 3.41e-20
C734 adder_4_2/adder_3_0/G1 A16 1.1e-19
C735 B12 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 3.81e-20
C736 SUB adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 1.39e-20
C737 adder_4_2/adder_3_0/G1 A13 9.55e-19
C738 S11 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_145_75# 1.39e-20
C739 adder_4_1/adder_3_0/P1 adder_4_2/adder_3_0/G2 5.87e-21
C740 adder_4_2/adder_3_0/P3 B15 2.06e-19
C741 adder_4_2/adder_3_0/P3 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 1.33e-20
C742 adder_4_3/CI adder_4_2/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# 6.93e-21
C743 S3 S4 -2e-23
C744 A15 adder_4_2/adder_3_0/G1 8.1e-20
C745 A5 adder_4_0/VDD 7.39e-21
C746 adder_4_2/CI B11 7.44e-19
C747 SUB S2 3.33e-22
C748 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# B15 4.06e-20
C749 SUB adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 1.17e-20
C750 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# B16 3.81e-20
C751 adder_4_1/adder_3_0/G2 adder_4_0/adder_3_0/P2 6.64e-21
C752 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# B8 2.14e-19
C753 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# S2 2.19e-20
C754 adder_4_0/VDD A7 2.34e-19
C755 B14 adder_4_2/adder_3_0/G2 6.51e-20
C756 adder_4_2/CI adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 3.7e-20
C757 S9 adder_4_3/adder_3_0/P3 1.67e-20
C758 A5 B6 1.11e-34
C759 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B B6 4.05e-19
C760 A8 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 6.43e-20
C761 B14 adder_4_3/VDD 5.55e-32
C762 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# CI 1.52e-20
C763 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B B15 1.18e-19
C764 adder_4_3/VDD adder_4_2/adder_3_0/P2 8.38e-19
C765 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 4.28e-21
C766 adder_4_2/CI adder_4_2/VDD 0.0264f
C767 adder_4_0/adder_3_0/G1 A5 9.55e-19
C768 adder_4_2/CI adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.433f
C769 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B B8 1.66e-19
C770 adder_4_1/adder_3_0/G1 A9 9.55e-19
C771 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# adder_4_1/CI 1.39e-35
C772 adder_4_1/VDD adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 4.75e-20
C773 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# A11 2.32e-20
C774 adder_4_1/adder_3_0/G3 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 2.84e-32
C775 adder_4_1/adder_3_0/P3 B12 5.72e-19
C776 adder_4_0/adder_3_0/G1 A7 8.1e-20
C777 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B A8 1.39e-19
C778 A14 adder_4_2/adder_3_0/P2 1.62e-19
C779 B16 adder_4_3/adder_3_0/G1 -6.94e-36
C780 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_4_3/CI 4.64e-20
C781 B8 adder_4_0/adder_2_0/G4 1.47e-21
C782 adder_4_3/CI adder_4_2/adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 4.91e-21
C783 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# S12 2.71e-19
C784 CI adder_4_1/adder_3_0/G1 0.0031f
C785 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# B8 3.81e-20
C786 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_4_1/CI 2.08e-19
C787 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_4_1/VDD 1.51e-19
C788 S3 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 5.56e-20
C789 B13 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 4.08e-21
C790 B9 adder_4_1/adder_3_0/G1 5.49e-20
C791 adder_4_1/adder_3_0/P3 adder_4_0/adder_3_0/P3 1.88e-19
C792 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# A8 3.19e-20
C793 B11 S5 8.93e-20
C794 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_2/adder_3_0/P1 4.66e-20
C795 SUB B12 0.00215f
C796 adder_4_1/CI adder_4_0/adder_2_0/G4 1.64e-21
C797 A7 adder_4_0/adder_3_0/G3 7.8e-20
C798 S5 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 6.6e-21
C799 SUB adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 3.41e-20
C800 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_4_1/VDD 2.78e-20
C801 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_4_1/CI 4.64e-20
C802 SUB adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 1.01e-20
C803 adder_4_3/adder_3_0/G2 B15 1.39e-35
C804 adder_4_1/adder_2_0/G4 adder_4_1/CI 3.53e-20
C805 adder_4_2/VDD S5 8.75e-19
C806 B16 adder_4_2/VDD 6.98e-19
C807 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 7.91e-21
C808 adder_4_1/adder_3_0/P3 A11 2.29e-19
C809 adder_4_2/adder_3_0/P2 B15 3.03e-19
C810 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# A12 6.43e-20
C811 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_4_2/adder_3_0/P2 2.53e-19
C812 SUB adder_4_0/adder_3_0/P3 1.14e-31
C813 SUB adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# 1.39e-20
C814 adder_4_1/adder_3_0/P3 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 3.3e-19
C815 adder_4_3/VDD adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 2.78e-20
C816 SUB B7 0.00112f
C817 B16 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 3.74e-19
C818 B8 adder_4_0/adder_3_0/P1 3.59e-19
C819 B6 CI 8.69e-19
C820 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B B8 3.74e-19
C821 A8 adder_4_0/adder_3_0/P1 2.81e-19
C822 adder_4_2/CI adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 2.46e-19
C823 B12 adder_4_2/CI 0.279f
C824 SUB adder_4_2/adder_3_0/G1 6.38e-21
C825 A8 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 1.4e-20
C826 SUB A11 8.93e-19
C827 A14 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 1.76e-20
C828 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_4_2/adder_3_0/G3 2.84e-32
C829 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 1.75e-20
C830 adder_4_2/adder_3_0/P3 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 1.97e-20
C831 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 5.8e-21
C832 adder_4_3/adder_3_0/P4 S12 2.69e-20
C833 adder_4_1/VDD adder_4_0/adder_3_0/P1 0.00122f
C834 adder_4_1/CI adder_4_0/adder_3_0/P1 4.71e-19
C835 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 7.69e-21
C836 S3 adder_4_1/adder_3_0/P4 2.35e-20
C837 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# B8 3.81e-20
C838 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_145_75# S3 1.39e-20
C839 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# B14 2.01e-20
C840 adder_4_1/adder_3_0/P2 B11 3.03e-19
C841 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_4_1/CI 5.9e-20
C842 adder_4_1/VDD adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 1.01e-19
C843 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# A8 3.19e-20
C844 B8 adder_4_0/adder_3_0/P2 4.43e-19
C845 S1 A7 1.1e-19
C846 B16 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 8.75e-20
C847 A16 S10 1.69e-19
C848 S1 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 5.99e-21
C849 A6 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 3.9e-19
C850 A6 adder_4_0/adder_3_0/P3 4.46e-20
C851 A8 adder_4_0/adder_3_0/P2 3.39e-19
C852 S8 A12 3.33e-19
C853 adder_4_0/adder_3_0/G2 B6 6.51e-20
C854 adder_4_1/adder_3_0/P2 adder_4_2/VDD 8.38e-19
C855 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_4_1/CI 4.64e-20
C856 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_4_1/VDD 5.65e-20
C857 S2 adder_4_1/adder_2_0/G4 1.98e-20
C858 A15 S10 3.71e-20
C859 B12 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 8.75e-20
C860 adder_4_1/VDD adder_4_0/adder_3_0/P2 8.38e-19
C861 adder_4_1/CI adder_4_0/adder_3_0/P2 6.08e-19
C862 adder_4_1/adder_3_0/G3 adder_4_1/CI 9.03e-20
C863 SUB adder_4_2/adder_2_0/G4 4.83e-20
C864 adder_4_1/adder_3_0/P1 B11 2.28e-19
C865 adder_4_2/CI A11 0.00338f
C866 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# B15 2.7e-20
C867 adder_4_2/adder_3_0/P2 adder_4_3/adder_3_0/P1 0.00296f
C868 adder_4_2/adder_3_0/P2 adder_4_1/CI 4.97e-20
C869 B12 S5 2.42e-19
C870 adder_4_1/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# adder_4_2/CI 3.27e-22
C871 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_0/adder_3_0/P1 4.66e-20
C872 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_4_3/CI 3.7e-20
C873 B11 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 1.18e-19
C874 adder_4_1/adder_3_0/P1 adder_4_2/VDD 0.00122f
C875 adder_4_1/adder_3_0/G3 B11 9.04e-20
C876 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 6.83e-22
C877 B16 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.00191f
C878 adder_4_1/CI adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 2.46e-19
C879 adder_4_2/adder_3_0/P2 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 5.27e-22
C880 B10 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 2.06e-22
C881 SUB A16 0.00154f
C882 adder_4_2/VDD adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 1.51e-19
C883 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_4_1/CI 2.04e-20
C884 SUB A13 1.99e-19
C885 adder_4_1/adder_3_0/G3 adder_4_2/VDD 5.85e-20
C886 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 3.19e-22
C887 B14 adder_4_2/VDD 2.46e-19
C888 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 3.22e-19
C889 adder_4_2/CI adder_4_2/adder_2_0/G4 3.53e-20
C890 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_4_0/adder_3_0/P2 2.19e-20
C891 S1 adder_4_1/adder_3_0/P4 1.83e-20
C892 SUB A15 8.93e-19
C893 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B A5 3.79e-20
C894 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 3.19e-22
C895 B12 adder_4_1/adder_2_0/G4 1.47e-21
C896 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 5e-21
C897 B10 A9 1.11e-34
C898 adder_4_2/adder_3_0/P2 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 3.15e-20
C899 B7 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 1.18e-19
C900 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# A12 4.77e-20
C901 B8 adder_4_1/adder_3_0/G1 -6.94e-36
C902 adder_4_0/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# B8 2.93e-22
C903 B16 adder_4_2/adder_3_0/G1 1.31e-19
C904 B14 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 2.79e-20
C905 S5 A11 1.1e-19
C906 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# B6 2.06e-22
C907 adder_4_2/adder_3_0/G3 adder_4_3/CI 1.54e-19
C908 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# 1.42e-19
C909 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B A7 4.82e-19
C910 A8 adder_4_1/adder_3_0/G1 -1.39e-35
C911 adder_4_3/VDD adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# -5.68e-32
C912 adder_4_2/CI adder_4_1/adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 4.91e-21
C913 adder_4_3/CI adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 1.39e-35
C914 adder_4_0/adder_2_0/sky130_fd_sc_hd__and4_1_0/X B8 3.37e-21
C915 adder_4_2/adder_3_0/P4 adder_4_2/CI 3.66e-20
C916 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_47# adder_4_1/CI 8.76e-20
C917 B12 adder_4_1/adder_3_0/P2 4.43e-19
C918 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_384_47# adder_4_1/adder_3_0/G2 4.9e-21
C919 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# B7 2.7e-20
C920 adder_4_2/adder_3_0/P1 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 6.6e-21
C921 adder_4_3/adder_3_0/G3 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 3.18e-20
C922 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# A12 4.77e-20
C923 adder_4_2/adder_3_0/P1 adder_4_3/adder_3_0/P2 1.07e-21
C924 B10 B9 -4.44e-34
C925 adder_4_1/VDD adder_4_1/adder_3_0/G1 2.84e-32
C926 adder_4_0/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# adder_4_1/CI 3.27e-22
C927 A16 adder_4_2/CI 5.12e-19
C928 adder_4_2/CI A13 3.01e-20
C929 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# S9 6.6e-21
C930 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_4_1/CI 1.52e-20
C931 adder_4_1/adder_3_0/P3 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 2.47e-20
C932 S4 adder_4_1/adder_3_0/P4 2.69e-20
C933 adder_4_2/adder_3_0/P1 adder_4_3/CI 4.71e-19
C934 adder_4_0/VDD B8 6.98e-19
C935 A15 adder_4_2/CI 2.75e-19
C936 adder_4_0/adder_2_0/sky130_fd_sc_hd__and4_1_0/X adder_4_1/CI 3.77e-21
C937 adder_4_1/adder_3_0/P2 adder_4_0/adder_3_0/P3 2.36e-20
C938 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_4_3/CI 4.64e-20
C939 A10 adder_4_1/adder_3_0/G2 5.72e-20
C940 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# B8 8.75e-20
C941 adder_4_0/VDD A8 6.31e-20
C942 B11 adder_4_1/adder_3_0/G1 9.39e-20
C943 B16 adder_4_2/adder_2_0/G4 1.47e-21
C944 adder_4_2/adder_2_0/G4 S5 1.75e-20
C945 B9 A12 5.55e-35
C946 SUB adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 1.76e-20
C947 B12 adder_4_1/adder_3_0/P1 3.59e-19
C948 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_4_0/adder_3_0/P1 6.6e-21
C949 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_47# CI 8.76e-20
C950 SUB S10 3.33e-22
C951 B10 adder_4_1/adder_3_0/G2 6.51e-20
C952 S6 A12 1.69e-19
C953 SUB adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 1.39e-20
C954 adder_4_3/VDD adder_4_2/adder_3_0/G3 5.85e-20
C955 adder_4_0/VDD adder_4_1/CI 0.00644f
C956 adder_4_0/adder_3_0/G1 B8 1.31e-19
C957 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# A12 3.71e-19
C958 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# adder_4_3/CI 2.04e-20
C959 A16 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 4.77e-20
C960 adder_4_2/VDD adder_4_1/adder_3_0/G1 5.65e-20
C961 B12 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 1.66e-19
C962 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_4_3/adder_3_0/P3 1.97e-20
C963 adder_4_1/adder_3_0/P2 A11 1.97e-19
C964 B7 adder_4_0/adder_3_0/P1 2.28e-19
C965 adder_4_3/VDD adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 4.75e-20
C966 adder_4_0/adder_3_0/G1 A8 1.1e-19
C967 A10 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 3.9e-19
C968 adder_4_2/CI adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 4.64e-20
C969 B12 adder_4_1/adder_3_0/G3 1.27e-19
C970 A16 S12 3.33e-19
C971 adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 0 0.00137f
C972 adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 0 0.255f
C973 A2 0 0.553f
C974 B2 0 0.632f
C975 adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 0 0.00137f
C976 adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 0 0.255f
C977 A1 0 0.469f
C978 B1 0 0.496f
C979 adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0 0.00137f
C980 adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 0 0.255f
C981 B4 0 1.05f
C982 A4 0 0.714f
C983 adder_4_0/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 0 0.177f
C984 B3 0 0.683f
C985 A3 0 0.729f
C986 adder_4_0/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 0 0.177f
C987 adder_4_0/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 0 0.177f
C988 adder_4_0/adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# 0 0.177f
C989 adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 0 0.00137f
C990 adder_4_0/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 0 0.255f
C991 S3 0 0.226f
C992 adder_4_0/adder_3_0/P3 0 1.49f
C993 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 0 0.00137f
C994 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 0 0.255f
C995 S2 0 0.212f
C996 adder_4_0/adder_3_0/P2 0 1.26f
C997 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 0 0.486f
C998 adder_4_0/VDD 0 17.4f
C999 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 0 0.00137f
C1000 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 0 0.255f
C1001 S1 0 0.353f
C1002 adder_4_0/adder_3_0/P1 0 1.11f
C1003 CI 0 2.13f
C1004 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0 0.00137f
C1005 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 0 0.255f
C1006 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 0 0.336f
C1007 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0 1.53f
C1008 adder_4_0/adder_3_0/G3 0 0.718f
C1009 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 0 0.0348f
C1010 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0 0.147f
C1011 adder_4_0/adder_3_0/G2 0 0.642f
C1012 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 0 0.0348f
C1013 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 0 0.147f
C1014 adder_4_0/adder_3_0/G1 0 0.527f
C1015 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# 0 0.0348f
C1016 adder_4_0/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 0 0.147f
C1017 S4 0 0.343f
C1018 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 0 0.00137f
C1019 adder_4_0/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 0 0.255f
C1020 adder_4_0/adder_2_0/sky130_fd_sc_hd__and4_1_0/X 0 0.154f
C1021 adder_4_0/adder_3_0/P4 0 1.62f
C1022 adder_4_0/adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 0 0.175f
C1023 adder_4_0/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# 0 0.0348f
C1024 adder_4_0/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# 0 0.147f
C1025 adder_4_0/adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 0 0.168f
C1026 adder_4_0/adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 0 0.129f
C1027 adder_4_0/adder_2_0/G4 0 0.596f
C1028 adder_4_0/adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 0 0.0348f
C1029 adder_4_0/adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0 0.147f
C1030 adder_4_0/adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 0 0.223f
C1031 adder_4_0/adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 0 0.0348f
C1032 adder_4_0/adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 0 0.147f
C1033 adder_4_0/adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# 0 0.0348f
C1034 adder_4_0/adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 0 0.147f
C1035 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 0 0.00137f
C1036 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 0 0.255f
C1037 A14 0 0.55f
C1038 B14 0 0.627f
C1039 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 0 0.00137f
C1040 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 0 0.255f
C1041 A13 0 0.467f
C1042 B13 0 0.491f
C1043 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0 0.00137f
C1044 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 0 0.255f
C1045 B16 0 1.05f
C1046 A16 0 0.714f
C1047 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 0 0.177f
C1048 B15 0 0.683f
C1049 A15 0 0.729f
C1050 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 0 0.177f
C1051 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 0 0.177f
C1052 adder_4_3/adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# 0 0.177f
C1053 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 0 0.00137f
C1054 adder_4_3/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 0 0.255f
C1055 S15 0 0.233f
C1056 adder_4_3/adder_3_0/P3 0 1.49f
C1057 adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 0 0.00137f
C1058 adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 0 0.255f
C1059 SUB 0 38.5f
C1060 S14 0 0.212f
C1061 adder_4_3/adder_3_0/P2 0 1.26f
C1062 adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 0 0.486f
C1063 adder_4_3/VDD 0 17.4f
C1064 adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 0 0.00137f
C1065 adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 0 0.255f
C1066 S13 0 0.353f
C1067 adder_4_3/adder_3_0/P1 0 1.11f
C1068 adder_4_3/CI 0 2.22f
C1069 adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0 0.00137f
C1070 adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 0 0.255f
C1071 adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 0 0.336f
C1072 adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0 1.53f
C1073 adder_4_3/adder_3_0/G3 0 0.718f
C1074 adder_4_3/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 0 0.0348f
C1075 adder_4_3/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0 0.147f
C1076 adder_4_3/adder_3_0/G2 0 0.642f
C1077 adder_4_3/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 0 0.0348f
C1078 adder_4_3/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 0 0.147f
C1079 adder_4_3/adder_3_0/G1 0 0.527f
C1080 adder_4_3/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# 0 0.0348f
C1081 adder_4_3/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 0 0.147f
C1082 S16 0 0.344f
C1083 adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 0 0.00137f
C1084 adder_4_3/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 0 0.255f
C1085 adder_4_3/adder_2_0/sky130_fd_sc_hd__and4_1_0/X 0 0.154f
C1086 adder_4_3/adder_3_0/P4 0 1.62f
C1087 adder_4_3/adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 0 0.175f
C1088 CO 0 0.959f
C1089 adder_4_3/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# 0 0.0348f
C1090 adder_4_3/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# 0 0.147f
C1091 adder_4_3/adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 0 0.168f
C1092 adder_4_3/adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 0 0.129f
C1093 adder_4_3/adder_2_0/G4 0 0.596f
C1094 adder_4_3/adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 0 0.0348f
C1095 adder_4_3/adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0 0.147f
C1096 adder_4_3/adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 0 0.223f
C1097 adder_4_3/adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 0 0.0348f
C1098 adder_4_3/adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 0 0.147f
C1099 adder_4_3/adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# 0 0.0348f
C1100 adder_4_3/adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 0 0.147f
C1101 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 0 0.00137f
C1102 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 0 0.255f
C1103 A10 0 0.55f
C1104 B10 0 0.627f
C1105 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 0 0.00137f
C1106 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 0 0.255f
C1107 A9 0 0.467f
C1108 B9 0 0.491f
C1109 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0 0.00137f
C1110 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 0 0.255f
C1111 B12 0 1.05f
C1112 A12 0 0.714f
C1113 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 0 0.177f
C1114 B11 0 0.683f
C1115 A11 0 0.729f
C1116 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 0 0.177f
C1117 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 0 0.177f
C1118 adder_4_2/adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# 0 0.177f
C1119 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 0 0.00137f
C1120 adder_4_2/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 0 0.255f
C1121 S11 0 0.226f
C1122 adder_4_2/adder_3_0/P3 0 1.49f
C1123 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 0 0.00137f
C1124 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 0 0.255f
C1125 S10 0 0.212f
C1126 adder_4_2/adder_3_0/P2 0 1.26f
C1127 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 0 0.486f
C1128 adder_4_2/VDD 0 17.4f
C1129 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 0 0.00137f
C1130 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 0 0.255f
C1131 S9 0 0.353f
C1132 adder_4_2/adder_3_0/P1 0 1.11f
C1133 adder_4_2/CI 0 2.23f
C1134 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0 0.00137f
C1135 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 0 0.255f
C1136 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 0 0.336f
C1137 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0 1.53f
C1138 adder_4_2/adder_3_0/G3 0 0.718f
C1139 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 0 0.0348f
C1140 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0 0.147f
C1141 adder_4_2/adder_3_0/G2 0 0.642f
C1142 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 0 0.0348f
C1143 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 0 0.147f
C1144 adder_4_2/adder_3_0/G1 0 0.527f
C1145 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# 0 0.0348f
C1146 adder_4_2/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 0 0.147f
C1147 S12 0 0.343f
C1148 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 0 0.00137f
C1149 adder_4_2/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 0 0.255f
C1150 adder_4_2/adder_2_0/sky130_fd_sc_hd__and4_1_0/X 0 0.154f
C1151 adder_4_2/adder_3_0/P4 0 1.62f
C1152 adder_4_2/adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 0 0.175f
C1153 adder_4_2/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# 0 0.0348f
C1154 adder_4_2/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# 0 0.147f
C1155 adder_4_2/adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 0 0.168f
C1156 adder_4_2/adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 0 0.129f
C1157 adder_4_2/adder_2_0/G4 0 0.596f
C1158 adder_4_2/adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 0 0.0348f
C1159 adder_4_2/adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0 0.147f
C1160 adder_4_2/adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 0 0.223f
C1161 adder_4_2/adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 0 0.0348f
C1162 adder_4_2/adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 0 0.147f
C1163 adder_4_2/adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# 0 0.0348f
C1164 adder_4_2/adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 0 0.147f
C1165 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 0 0.00137f
C1166 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 0 0.255f
C1167 A6 0 0.55f
C1168 B6 0 0.627f
C1169 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 0 0.00137f
C1170 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 0 0.255f
C1171 A5 0 0.467f
C1172 B5 0 0.491f
C1173 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0 0.00137f
C1174 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 0 0.255f
C1175 B8 0 1.05f
C1176 A8 0 0.714f
C1177 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 0 0.177f
C1178 B7 0 0.683f
C1179 A7 0 0.729f
C1180 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 0 0.177f
C1181 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 0 0.177f
C1182 adder_4_1/adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# 0 0.177f
C1183 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 0 0.00137f
C1184 adder_4_1/adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 0 0.255f
C1185 S7 0 0.226f
C1186 adder_4_1/adder_3_0/P3 0 1.49f
C1187 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 0 0.00137f
C1188 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 0 0.255f
C1189 S6 0 0.212f
C1190 adder_4_1/adder_3_0/P2 0 1.26f
C1191 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 0 0.486f
C1192 adder_4_1/VDD 0 17.4f
C1193 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 0 0.00137f
C1194 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 0 0.255f
C1195 S5 0 0.353f
C1196 adder_4_1/adder_3_0/P1 0 1.11f
C1197 adder_4_1/CI 0 2.22f
C1198 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0 0.00137f
C1199 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 0 0.255f
C1200 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 0 0.336f
C1201 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0 1.53f
C1202 adder_4_1/adder_3_0/G3 0 0.718f
C1203 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 0 0.0348f
C1204 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0 0.147f
C1205 adder_4_1/adder_3_0/G2 0 0.642f
C1206 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 0 0.0348f
C1207 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 0 0.147f
C1208 adder_4_1/adder_3_0/G1 0 0.527f
C1209 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# 0 0.0348f
C1210 adder_4_1/adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 0 0.147f
C1211 S8 0 0.343f
C1212 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 0 0.00137f
C1213 adder_4_1/adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 0 0.255f
C1214 adder_4_1/adder_2_0/sky130_fd_sc_hd__and4_1_0/X 0 0.154f
C1215 adder_4_1/adder_3_0/P4 0 1.62f
C1216 adder_4_1/adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 0 0.175f
C1217 adder_4_1/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# 0 0.0348f
C1218 adder_4_1/adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# 0 0.147f
C1219 adder_4_1/adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 0 0.168f
C1220 adder_4_1/adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 0 0.129f
C1221 adder_4_1/adder_2_0/G4 0 0.596f
C1222 adder_4_1/adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 0 0.0348f
C1223 adder_4_1/adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0 0.147f
C1224 adder_4_1/adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 0 0.223f
C1225 adder_4_1/adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 0 0.0348f
C1226 adder_4_1/adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 0 0.147f
C1227 adder_4_1/adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# 0 0.0348f
C1228 adder_4_1/adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 0 0.147f
.ends

