magic
tech sky130A
magscale 1 2
timestamp 1704906721
<< nwell >>
rect 570 264 596 585
rect 1212 264 1231 585
rect 1850 580 2110 585
rect 1850 264 1860 580
rect 2736 264 2758 585
rect 3461 264 3484 585
rect 4194 264 4220 585
<< pwell >>
rect 537 51 634 206
rect 1170 51 1269 206
rect 1810 51 1905 200
rect 1971 51 2078 198
rect 2701 51 2804 205
rect 3423 51 3532 206
rect 4152 51 4262 206
<< locali >>
rect 542 530 575 564
rect 610 530 636 564
rect 1171 530 1205 564
rect 1240 530 1269 564
rect 1803 530 1840 564
rect 1875 530 1898 564
rect 1973 530 2010 564
rect 2045 530 2069 564
rect 2704 530 2731 564
rect 2766 530 2798 564
rect 3423 530 3461 564
rect 3496 530 3525 564
rect 4153 530 4186 564
rect 4221 530 4255 564
rect 665 460 699 462
rect 660 430 699 460
rect 690 428 699 430
rect 1300 428 1334 462
rect 690 425 695 428
rect 30 340 64 345
rect 657 325 691 326
rect 542 -14 570 20
rect 605 -14 632 20
rect 1175 -14 1205 20
rect 1240 -14 1268 20
rect 1805 -14 1840 20
rect 1875 -14 1899 20
rect 1984 -14 2010 20
rect 2045 -14 2068 20
rect 2697 -14 2731 20
rect 2766 -14 2793 20
rect 3424 -14 3456 20
rect 3491 -14 3528 20
rect 4159 -14 4186 20
rect 4221 -14 4255 20
<< viali >>
rect 575 530 610 564
rect 1205 530 1240 564
rect 1840 530 1875 564
rect 2010 530 2045 564
rect 2731 530 2766 564
rect 3461 530 3496 564
rect 4186 530 4221 564
rect 655 395 690 430
rect 25 305 60 340
rect 2631 310 2665 344
rect 3356 310 3390 344
rect 4086 310 4120 344
rect 4816 310 4850 344
rect 217 218 251 252
rect 345 218 379 252
rect 473 218 507 252
rect 852 218 886 252
rect 980 218 1014 252
rect 1108 218 1142 252
rect 1487 218 1521 252
rect 1615 218 1649 252
rect 1743 218 1777 252
rect 2149 218 2183 252
rect 2266 218 2300 252
rect 2874 218 2908 252
rect 2991 218 3025 252
rect 3604 218 3638 252
rect 3721 218 3755 252
rect 4334 218 4368 252
rect 4451 218 4485 252
rect 1295 120 1330 155
rect 570 -14 605 20
rect 1205 -14 1240 20
rect 1840 -14 1875 20
rect 2010 -14 2045 20
rect 2731 -14 2766 20
rect 3456 -14 3491 20
rect 4186 -14 4221 20
<< metal1 >>
rect 480 590 520 595
rect 541 564 631 595
rect 541 530 575 564
rect 610 530 631 564
rect 541 499 631 530
rect 1178 564 1270 595
rect 1178 530 1205 564
rect 1240 530 1270 564
rect 1178 499 1270 530
rect 1810 564 1898 595
rect 1810 530 1840 564
rect 1875 530 1898 564
rect 1810 499 1898 530
rect 1982 564 2071 595
rect 1982 530 2010 564
rect 2045 530 2071 564
rect 1982 499 2071 530
rect 2699 564 2793 595
rect 2699 530 2731 564
rect 2766 530 2793 564
rect 2699 499 2793 530
rect 3428 564 3523 595
rect 3428 530 3461 564
rect 3496 530 3523 564
rect 3428 499 3523 530
rect 4158 564 4255 595
rect 4158 530 4186 564
rect 4221 530 4255 564
rect 4158 499 4255 530
rect 635 445 715 455
rect 635 385 645 445
rect 705 385 715 445
rect 635 375 715 385
rect 2611 355 2691 365
rect 10 340 70 350
rect 10 305 25 340
rect 60 310 2550 340
rect 60 305 70 310
rect 10 290 70 305
rect 190 270 270 280
rect 190 210 200 270
rect 260 210 270 270
rect 190 200 270 210
rect 315 270 395 280
rect 315 210 325 270
rect 385 210 395 270
rect 315 200 395 210
rect 455 270 535 280
rect 980 275 1010 310
rect 455 210 465 270
rect 525 210 535 270
rect 455 200 535 210
rect 825 265 905 275
rect 825 205 835 265
rect 895 205 905 265
rect 825 195 905 205
rect 955 265 1035 275
rect 955 205 965 265
rect 1025 205 1035 265
rect 955 195 1035 205
rect 1085 265 1165 275
rect 1085 205 1095 265
rect 1155 205 1165 265
rect 1085 195 1165 205
rect 1460 265 1540 275
rect 1460 205 1470 265
rect 1530 205 1540 265
rect 1460 195 1540 205
rect 1585 265 1665 275
rect 1585 205 1595 265
rect 1655 205 1665 265
rect 1585 195 1665 205
rect 1725 265 1805 275
rect 1725 205 1735 265
rect 1795 205 1805 265
rect 1725 195 1805 205
rect 2126 260 2206 270
rect 2126 200 2136 260
rect 2196 200 2206 260
rect 2126 190 2206 200
rect 2246 265 2326 275
rect 2246 205 2256 265
rect 2316 205 2326 265
rect 2520 250 2550 310
rect 2611 295 2621 355
rect 2681 295 2691 355
rect 2611 285 2691 295
rect 3336 350 3416 360
rect 3336 295 3346 350
rect 3406 295 3416 350
rect 3336 285 3416 295
rect 4066 355 4146 365
rect 4066 295 4076 355
rect 4136 295 4146 355
rect 4066 285 4146 295
rect 4796 355 4876 365
rect 4796 300 4806 355
rect 4866 300 4876 355
rect 4796 290 4876 300
rect 2851 270 2931 280
rect 2851 250 2861 270
rect 2520 220 2861 250
rect 2246 195 2326 205
rect 2851 210 2861 220
rect 2921 210 2931 270
rect 3581 265 3661 275
rect 2851 200 2931 210
rect 2966 255 3046 265
rect 2966 195 2976 255
rect 3036 195 3046 255
rect 3581 205 3591 265
rect 3651 205 3661 265
rect 3581 195 3661 205
rect 3696 265 3776 275
rect 3696 205 3706 265
rect 3766 205 3776 265
rect 3696 195 3776 205
rect 4311 265 4391 275
rect 4311 205 4321 265
rect 4381 205 4391 265
rect 4311 195 4391 205
rect 4426 265 4506 275
rect 4426 205 4436 265
rect 4496 205 4506 265
rect 4426 195 4506 205
rect 2966 185 3046 195
rect 1280 155 1340 165
rect 4335 155 4365 195
rect 1280 120 1295 155
rect 1330 125 4365 155
rect 1330 120 1340 125
rect 1280 105 1340 120
rect 539 20 636 51
rect 539 -14 570 20
rect 605 -14 636 20
rect 539 -45 636 -14
rect 1167 20 1269 51
rect 1167 -14 1205 20
rect 1240 -14 1269 20
rect 1167 -45 1269 -14
rect 1810 20 1902 51
rect 1810 -14 1840 20
rect 1875 -14 1902 20
rect 1810 -45 1902 -14
rect 1978 20 2068 51
rect 1978 -14 2010 20
rect 2045 -14 2068 20
rect 1978 -45 2068 -14
rect 2704 20 2794 51
rect 2704 -14 2731 20
rect 2766 -14 2794 20
rect 2704 -45 2794 -14
rect 3428 20 3524 51
rect 3428 -14 3456 20
rect 3491 -14 3524 20
rect 3428 -45 3524 -14
rect 4158 20 4255 51
rect 4158 -14 4186 20
rect 4221 -14 4255 20
rect 4158 -45 4255 -14
rect 450 -85 530 -75
rect 450 -145 460 -85
rect 520 -100 530 -85
rect 2245 -85 2325 -75
rect 2245 -100 2255 -85
rect 520 -130 2255 -100
rect 520 -145 530 -130
rect 450 -155 530 -145
rect 2245 -145 2255 -130
rect 2315 -145 2325 -85
rect 2245 -155 2325 -145
rect 1085 -170 1165 -160
rect 1085 -230 1095 -170
rect 1155 -185 1165 -170
rect 2965 -170 3045 -160
rect 2965 -185 2975 -170
rect 1155 -215 2975 -185
rect 1155 -230 1165 -215
rect 1085 -240 1165 -230
rect 2965 -230 2975 -215
rect 3035 -230 3045 -170
rect 2965 -240 3045 -230
rect 1720 -255 1800 -245
rect 1720 -315 1730 -255
rect 1790 -270 1800 -255
rect 3700 -255 3780 -245
rect 3700 -270 3710 -255
rect 1790 -300 3710 -270
rect 1790 -315 1800 -300
rect 1720 -325 1800 -315
rect 3700 -315 3710 -300
rect 3770 -315 3780 -255
rect 3700 -325 3780 -315
rect 325 -340 405 -330
rect 325 -400 335 -340
rect 395 -355 405 -340
rect 2125 -340 2205 -330
rect 2125 -355 2135 -340
rect 395 -385 2135 -355
rect 395 -400 405 -385
rect 325 -410 405 -400
rect 2125 -400 2135 -385
rect 2195 -400 2205 -340
rect 2125 -410 2205 -400
rect 630 -425 710 -415
rect 630 -485 640 -425
rect 700 -440 710 -425
rect 1590 -425 1670 -415
rect 1590 -440 1600 -425
rect 700 -470 1600 -440
rect 700 -485 710 -470
rect 630 -495 710 -485
rect 1590 -485 1600 -470
rect 1660 -440 1670 -425
rect 3580 -425 3660 -415
rect 3580 -440 3590 -425
rect 1660 -470 3590 -440
rect 1660 -485 1670 -470
rect 1590 -495 1670 -485
rect 3580 -485 3590 -470
rect 3650 -485 3660 -425
rect 3580 -495 3660 -485
<< via1 >>
rect 645 430 705 445
rect 645 395 655 430
rect 655 395 690 430
rect 690 395 705 430
rect 645 385 705 395
rect 200 252 260 270
rect 200 218 217 252
rect 217 218 251 252
rect 251 218 260 252
rect 200 210 260 218
rect 325 252 385 270
rect 325 218 345 252
rect 345 218 379 252
rect 379 218 385 252
rect 325 210 385 218
rect 465 252 525 270
rect 465 218 473 252
rect 473 218 507 252
rect 507 218 525 252
rect 465 210 525 218
rect 835 252 895 265
rect 835 218 852 252
rect 852 218 886 252
rect 886 218 895 252
rect 835 205 895 218
rect 965 252 1025 265
rect 965 218 980 252
rect 980 218 1014 252
rect 1014 218 1025 252
rect 965 205 1025 218
rect 1095 252 1155 265
rect 1095 218 1108 252
rect 1108 218 1142 252
rect 1142 218 1155 252
rect 1095 205 1155 218
rect 1470 252 1530 265
rect 1470 218 1487 252
rect 1487 218 1521 252
rect 1521 218 1530 252
rect 1470 205 1530 218
rect 1595 252 1655 265
rect 1595 218 1615 252
rect 1615 218 1649 252
rect 1649 218 1655 252
rect 1595 205 1655 218
rect 1735 252 1795 265
rect 1735 218 1743 252
rect 1743 218 1777 252
rect 1777 218 1795 252
rect 1735 205 1795 218
rect 2136 252 2196 260
rect 2136 218 2149 252
rect 2149 218 2183 252
rect 2183 218 2196 252
rect 2136 200 2196 218
rect 2256 252 2316 265
rect 2256 218 2266 252
rect 2266 218 2300 252
rect 2300 218 2316 252
rect 2256 205 2316 218
rect 2621 344 2681 355
rect 2621 310 2631 344
rect 2631 310 2665 344
rect 2665 310 2681 344
rect 2621 295 2681 310
rect 3346 344 3406 350
rect 3346 310 3356 344
rect 3356 310 3390 344
rect 3390 310 3406 344
rect 3346 295 3406 310
rect 4076 344 4136 355
rect 4076 310 4086 344
rect 4086 310 4120 344
rect 4120 310 4136 344
rect 4076 295 4136 310
rect 4806 344 4866 355
rect 4806 310 4816 344
rect 4816 310 4850 344
rect 4850 310 4866 344
rect 4806 300 4866 310
rect 2861 252 2921 270
rect 2861 218 2874 252
rect 2874 218 2908 252
rect 2908 218 2921 252
rect 2861 210 2921 218
rect 2976 252 3036 255
rect 2976 218 2991 252
rect 2991 218 3025 252
rect 3025 218 3036 252
rect 2976 195 3036 218
rect 3591 252 3651 265
rect 3591 218 3604 252
rect 3604 218 3638 252
rect 3638 218 3651 252
rect 3591 205 3651 218
rect 3706 252 3766 265
rect 3706 218 3721 252
rect 3721 218 3755 252
rect 3755 218 3766 252
rect 3706 205 3766 218
rect 4321 252 4381 265
rect 4321 218 4334 252
rect 4334 218 4368 252
rect 4368 218 4381 252
rect 4321 205 4381 218
rect 4436 252 4496 265
rect 4436 218 4451 252
rect 4451 218 4485 252
rect 4485 218 4496 252
rect 4436 205 4496 218
rect 460 -145 520 -85
rect 2255 -145 2315 -85
rect 1095 -230 1155 -170
rect 2975 -230 3035 -170
rect 1730 -315 1790 -255
rect 3710 -315 3770 -255
rect 335 -400 395 -340
rect 2135 -400 2195 -340
rect 640 -485 700 -425
rect 1600 -485 1660 -425
rect 3590 -485 3650 -425
<< metal2 >>
rect 635 445 715 455
rect 635 385 645 445
rect 705 385 715 445
rect 635 375 715 385
rect 190 270 270 280
rect 190 210 200 270
rect 260 210 270 270
rect 190 200 270 210
rect 315 270 395 280
rect 315 210 325 270
rect 385 210 395 270
rect 315 200 395 210
rect 455 270 535 280
rect 455 210 465 270
rect 525 210 535 270
rect 455 200 535 210
rect 350 -330 380 200
rect 475 -75 505 200
rect 450 -85 530 -75
rect 450 -145 460 -85
rect 520 -145 530 -85
rect 450 -155 530 -145
rect 325 -340 405 -330
rect 325 -400 335 -340
rect 395 -400 405 -340
rect 325 -410 405 -400
rect 655 -415 685 375
rect 2611 355 2691 365
rect 2611 295 2621 355
rect 2681 295 2691 355
rect 2611 285 2691 295
rect 3336 350 3416 360
rect 3336 295 3346 350
rect 3406 295 3416 350
rect 3336 285 3416 295
rect 4066 355 4146 365
rect 4066 295 4076 355
rect 4136 295 4146 355
rect 4066 285 4146 295
rect 4796 355 4876 365
rect 4796 300 4806 355
rect 4866 300 4876 355
rect 4796 290 4876 300
rect 825 265 905 275
rect 825 205 835 265
rect 895 205 905 265
rect 825 195 905 205
rect 955 265 1035 275
rect 955 205 965 265
rect 1025 205 1035 265
rect 955 195 1035 205
rect 1085 265 1165 275
rect 1085 205 1095 265
rect 1155 205 1165 265
rect 1085 195 1165 205
rect 1460 265 1540 275
rect 1460 205 1470 265
rect 1530 205 1540 265
rect 1460 195 1540 205
rect 1585 265 1665 275
rect 1585 205 1595 265
rect 1655 205 1665 265
rect 1585 195 1665 205
rect 1725 265 1805 275
rect 1725 205 1735 265
rect 1795 205 1805 265
rect 1110 -160 1140 195
rect 1085 -170 1165 -160
rect 1085 -230 1095 -170
rect 1155 -230 1165 -170
rect 1085 -240 1165 -230
rect 1615 -415 1645 195
rect 1725 194 1805 205
rect 2126 260 2206 270
rect 2126 200 2136 260
rect 2196 200 2206 260
rect 1745 -245 1775 194
rect 2126 190 2206 200
rect 2246 265 2326 275
rect 2246 205 2256 265
rect 2316 205 2326 265
rect 2246 195 2326 205
rect 2851 270 2931 280
rect 2851 210 2861 270
rect 2921 210 2931 270
rect 3581 265 3661 275
rect 2851 200 2931 210
rect 2966 255 3046 265
rect 2966 195 2976 255
rect 3036 195 3046 255
rect 3581 205 3591 265
rect 3651 205 3661 265
rect 3581 195 3661 205
rect 3696 265 3776 275
rect 3696 205 3706 265
rect 3766 205 3776 265
rect 3696 195 3776 205
rect 4311 265 4391 275
rect 4311 205 4321 265
rect 4381 205 4391 265
rect 4311 195 4391 205
rect 4426 265 4506 275
rect 4426 205 4436 265
rect 4496 205 4506 265
rect 4426 195 4506 205
rect 1720 -255 1800 -245
rect 1720 -315 1730 -255
rect 1790 -315 1800 -255
rect 1720 -325 1800 -315
rect 2150 -330 2180 190
rect 2270 -75 2300 195
rect 2966 185 3046 195
rect 2245 -85 2325 -75
rect 2245 -145 2255 -85
rect 2315 -145 2325 -85
rect 2245 -155 2325 -145
rect 2990 -160 3020 185
rect 2965 -170 3045 -160
rect 2965 -230 2975 -170
rect 3035 -230 3045 -170
rect 2965 -240 3045 -230
rect 2125 -340 2205 -330
rect 2125 -400 2135 -340
rect 2195 -400 2205 -340
rect 2125 -410 2205 -400
rect 3605 -415 3635 195
rect 3725 -245 3755 195
rect 3700 -255 3780 -245
rect 3700 -315 3710 -255
rect 3770 -315 3780 -255
rect 3700 -325 3780 -315
rect 630 -425 710 -415
rect 630 -485 640 -425
rect 700 -485 710 -425
rect 630 -495 710 -485
rect 1590 -425 1670 -415
rect 1590 -485 1600 -425
rect 1660 -485 1670 -425
rect 1590 -495 1670 -485
rect 3580 -425 3660 -415
rect 3580 -485 3590 -425
rect 3650 -485 3660 -425
rect 3580 -495 3660 -485
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_0
timestamp 1691611044
transform 1 0 -7 0 1 3
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_1
timestamp 1691611044
transform 1 0 628 0 1 3
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_2
timestamp 1691611044
transform 1 0 1263 0 1 3
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1691611044
transform 1 0 1896 0 1 3
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_0
timestamp 1691611044
transform 1 0 2064 0 1 3
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_1
timestamp 1691611044
transform 1 0 2789 0 1 3
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_2
timestamp 1691611044
transform 1 0 3519 0 1 3
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_3
timestamp 1691611044
transform 1 0 4249 0 1 3
box -38 -48 682 592
<< labels >>
flabel via1 490 240 490 240 1 FreeSans 128 0 0 0 P1
port 2 n
flabel via1 360 240 360 240 1 FreeSans 160 0 0 0 CI
port 1 n
flabel via1 1125 235 1125 235 1 FreeSans 240 0 0 0 P2
port 4 n
flabel via1 234 240 234 240 1 FreeSans 128 0 0 0 G1
port 3 n
flabel via1 870 240 870 240 1 FreeSans 160 0 0 0 G2
port 5 n
flabel via1 1760 245 1760 245 1 FreeSans 128 0 0 0 P3
port 6 n
flabel via1 1500 245 1500 245 1 FreeSans 128 0 0 0 G3
port 7 n
flabel metal1 s 555 35 555 35 1 FreeSans 160 0 0 0 GND
port 16 n
flabel viali s 595 550 595 550 1 FreeSans 160 0 0 0 VDD
port 15 n
flabel via1 3371 335 3371 335 1 FreeSans 128 0 0 0 S2
port 11 n
flabel via1 4101 335 4101 335 1 FreeSans 160 0 0 0 S3
port 12 n
flabel via1 4831 335 4831 335 1 FreeSans 160 0 0 0 S4
port 13 n
flabel via1 2646 335 2646 335 1 FreeSans 128 0 0 0 S1
port 10 n
flabel nwell s 1935 350 1935 350 1 FreeSans 240 0 0 0 VPB
port 17 n
flabel via1 4467 241 4467 241 1 FreeSans 64 0 0 0 P4
port 8 n
<< end >>
