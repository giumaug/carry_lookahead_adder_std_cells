ADDER_4

v1 CI GND pwl 0 0ps
v2 A4 GND pwl 0 0ps
v3 B4 GND pwl 0 0ps 1000ps 0 1050ps 1.8
v4 A3 GND pwl 0 0ps
v5 B3 GND pwl 0 0ps 1000ps 0 1050ps 1.8
v6 A2 GND pwl 0 0ps
v7 B2 GND pwl 0 0ps 1000ps 0 1050ps 1.8
v8 A1 GND pwl 0 0ps 1000ps 0 1050ps 1.8
v9 B1 GND pwl 0 0ps 1000ps 0 1050ps 1.8
v10 VDD GND pwl 0 1.8

Xadder_4_0 A1 B1 A2 B2 A3 B3 A4 B4 CI S1 S2 S3 S4 CO VDD GND adder_4

.measure tran tpdr TRIG v(B1) VAL=0.1 RISE=1 TARG v(co) VAL=1.7 RISE=1
*.measure tran tpdf TRIG v(B1) VAL=1.7 FALL=1 TARG v(co) VAL=0.1 FALL=1 CROSS=LAST


.lib /opt/open_pdks/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt
*.tran 10p 204800ps
*.options method=gear
*.tran 40ps 4000ps
*.save all

.control
tran 40ps 4000ps
options method=gear
let ret = v(co)[length(co)-1]
echo $&ret >> xxx.txt
.endc

.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X a_384_47# a_81_21# a_299_297#
X0 a_81_21# B1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0894 pd=0.925 as=0.229 ps=1.57 w=0.65 l=0.15
**devattr s=10270,288 d=3575,185
X1 a_299_297# B1 a_81_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.69 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5500,255
X2 VPWR a_81_21# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.69 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=10400,504
X3 VPWR A1 a_299_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.69 as=0.18 ps=1.69 w=1 l=0.15
**devattr s=5500,255 d=5600,256
X4 VGND a_81_21# X VNB sky130_fd_pr__nfet_01v8 ad=0.229 pd=1.57 as=0.169 ps=1.82 w=0.65 l=0.15
**devattr s=6760,364 d=10270,288
X5 VGND A2 a_384_47# VNB sky130_fd_pr__nfet_01v8 ad=0.229 pd=1.57 as=0.091 ps=0.93 w=0.65 l=0.15
**devattr s=3640,186 d=6890,366
X6 a_299_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.69 as=0.18 ps=1.69 w=1 l=0.15
**devattr s=5600,256 d=10600,506
X7 a_384_47# A1 a_81_21# VNB sky130_fd_pr__nfet_01v8 ad=0.091 pd=0.93 as=0.0894 ps=0.925 w=0.65 l=0.15
**devattr s=3575,185 d=3640,186
C0 B1 A1 0.0817f
C1 X a_81_21# 0.112f
C2 X VPB 0.0108f
C3 a_299_297# VGND 0.00772f
C4 VGND a_81_21# 0.173f
C5 VPWR A1 0.0209f
C6 VGND VPB 0.00713f
C7 VPWR A2 0.0201f
C8 X B1 3.04e-20
C9 a_299_297# a_81_21# 0.0821f
C10 a_299_297# VPB 0.0111f
C11 a_81_21# VPB 0.0593f
C12 VGND B1 0.0181f
C13 a_384_47# A1 0.00884f
C14 X VPWR 0.0847f
C15 VPWR VGND 0.0579f
C16 a_299_297# B1 0.00863f
C17 a_81_21# B1 0.148f
C18 B1 VPB 0.0387f
C19 a_299_297# VPWR 0.202f
C20 A1 A2 0.0921f
C21 VPWR a_81_21# 0.146f
C22 VPWR VPB 0.068f
C23 a_384_47# VGND 0.00366f
C24 a_299_297# a_384_47# 1.48e-19
C25 VPWR B1 0.0196f
C26 a_384_47# a_81_21# 0.00138f
C27 VGND A1 0.0786f
C28 VGND A2 0.0495f
C29 a_299_297# A1 0.0585f
C30 a_81_21# A1 0.0568f
C31 a_299_297# A2 0.0468f
C32 a_81_21# A2 7.47e-19
C33 A1 VPB 0.0264f
C34 X VGND 0.0512f
C35 A2 VPB 0.0373f
C36 a_384_47# VPWR 4.08e-19
C37 VGND VNB 0.364f
C38 VPWR VNB 0.286f
C39 X VNB 0.0945f
C40 A2 VNB 0.144f
C41 A1 VNB 0.0996f
C42 B1 VNB 0.109f
C43 VPB VNB 0.605f
C44 a_299_297# VNB 0.0348f
C45 a_81_21# VNB 0.147f
.ends

.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X a_109_47# a_197_47# a_303_47#
+ a_27_47#
X0 a_27_47# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.139 ps=0.987 w=0.42 l=0.15
**devattr s=3108,158 d=2352,140
X1 a_197_47# B a_109_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0798 pd=0.8 as=0.0609 ps=0.71 w=0.42 l=0.15
**devattr s=2436,142 d=3192,160
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.332 ps=2.35 w=1 l=0.15
**devattr s=12498,336 d=10400,504
X3 a_303_47# C a_197_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0798 ps=0.8 w=0.42 l=0.15
**devattr s=3192,160 d=2772,150
X4 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0662 pd=0.735 as=0.139 ps=0.987 w=0.42 l=0.15
**devattr s=4368,272 d=2940,154
X5 VPWR D a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.139 pd=0.987 as=0.0662 ps=0.735 w=0.42 l=0.15
**devattr s=2352,140 d=12498,336
X6 VGND D a_303_47# VNB sky130_fd_pr__nfet_01v8 ad=0.154 pd=1.04 as=0.0693 ps=0.75 w=0.42 l=0.15
**devattr s=2772,150 d=7851,266
X7 VPWR B a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.139 pd=0.987 as=0.0662 ps=0.735 w=0.42 l=0.15
**devattr s=2940,154 d=3108,158
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.238 ps=1.62 w=0.65 l=0.15
**devattr s=7851,266 d=6760,364
X9 a_109_47# A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.109 ps=1.36 w=0.42 l=0.15
**devattr s=4368,272 d=2436,142
C0 VPB a_27_47# 0.082f
C1 VGND A 0.0151f
C2 C a_109_47# 1.72e-20
C3 A a_27_47# 0.153f
C4 VGND a_27_47# 0.132f
C5 D VPWR 0.0207f
C6 VPB X 0.0111f
C7 D a_303_47# 0.00119f
C8 C D 0.18f
C9 X VGND 0.0903f
C10 VGND a_109_47# 0.00223f
C11 B VPWR 0.0231f
C12 B a_197_47# 0.00623f
C13 X a_27_47# 0.0754f
C14 a_109_47# a_27_47# 0.00578f
C15 VPWR a_197_47# 5.24e-19
C16 D VPB 0.0782f
C17 VPWR a_303_47# 4.83e-19
C18 C B 0.161f
C19 C VPWR 0.021f
C20 D VGND 0.0898f
C21 C a_197_47# 0.00123f
C22 C a_303_47# 0.00527f
C23 D a_27_47# 0.107f
C24 B VPB 0.0643f
C25 VPB VPWR 0.077f
C26 B A 0.0839f
C27 A VPWR 0.044f
C28 B VGND 0.0453f
C29 VGND VPWR 0.0662f
C30 D X 0.00746f
C31 C VPB 0.0609f
C32 VGND a_197_47# 0.00387f
C33 VGND a_303_47# 0.00381f
C34 B a_27_47# 0.13f
C35 VPWR a_27_47# 0.326f
C36 a_197_47# a_27_47# 0.00167f
C37 a_303_47# a_27_47# 0.00119f
C38 C VGND 0.0408f
C39 VPB A 0.0907f
C40 C a_27_47# 0.0516f
C41 X VPWR 0.0945f
C42 B a_109_47# 0.00153f
C43 VPWR a_109_47# 4.66e-19
C44 VPB VGND 0.00852f
C45 VGND VNB 0.393f
C46 X VNB 0.0933f
C47 VPWR VNB 0.335f
C48 D VNB 0.13f
C49 C VNB 0.11f
C50 B VNB 0.112f
C51 A VNB 0.221f
C52 VPB VNB 0.693f
C53 a_27_47# VNB 0.175f
.ends

.subckt adder_2 CI P1 G1 P2 G2 P3 G3 P4 G4 CO sky130_fd_sc_hd__a21o_1_0/a_81_21# sky130_fd_sc_hd__and4_1_0/a_27_47#
+ sky130_fd_sc_hd__a21o_1_0/a_384_47# sky130_fd_sc_hd__a21o_1_1/X sky130_fd_sc_hd__a21o_1_1/a_81_21#
+ sky130_fd_sc_hd__a21o_1_0/a_299_297# VPB sky130_fd_sc_hd__a21o_1_1/a_299_297# sky130_fd_sc_hd__a21o_1_1/a_384_47#
+ sky130_fd_sc_hd__a21o_1_2/a_299_297# sky130_fd_sc_hd__and4_1_0/a_109_47# sky130_fd_sc_hd__a21o_1_2/X
+ sky130_fd_sc_hd__a21o_1_0/X sky130_fd_sc_hd__and4_1_0/X sky130_fd_sc_hd__a21o_1_3/a_299_297#
+ sky130_fd_sc_hd__a21o_1_2/a_81_21# VNB sky130_fd_sc_hd__and4_1_0/a_197_47# sky130_fd_sc_hd__a21o_1_2/a_384_47#
+ sky130_fd_sc_hd__and4_1_0/a_303_47# sky130_fd_sc_hd__a21o_1_3/a_81_21# sky130_fd_sc_hd__a21o_1_3/a_384_47#
Xsky130_fd_sc_hd__a21o_1_0 G1 P2 G2 VNB VNB VPB VPB sky130_fd_sc_hd__a21o_1_0/X sky130_fd_sc_hd__a21o_1_0/a_384_47#
+ sky130_fd_sc_hd__a21o_1_0/a_81_21# sky130_fd_sc_hd__a21o_1_0/a_299_297# sky130_fd_sc_hd__a21o_1
Xsky130_fd_sc_hd__a21o_1_1 sky130_fd_sc_hd__a21o_1_0/X P3 G3 VNB VNB VPB VPB sky130_fd_sc_hd__a21o_1_1/X
+ sky130_fd_sc_hd__a21o_1_1/a_384_47# sky130_fd_sc_hd__a21o_1_1/a_81_21# sky130_fd_sc_hd__a21o_1_1/a_299_297#
+ sky130_fd_sc_hd__a21o_1
Xsky130_fd_sc_hd__a21o_1_2 sky130_fd_sc_hd__a21o_1_1/X P4 G4 VNB VNB VPB VPB sky130_fd_sc_hd__a21o_1_2/X
+ sky130_fd_sc_hd__a21o_1_2/a_384_47# sky130_fd_sc_hd__a21o_1_2/a_81_21# sky130_fd_sc_hd__a21o_1_2/a_299_297#
+ sky130_fd_sc_hd__a21o_1
Xsky130_fd_sc_hd__a21o_1_3 sky130_fd_sc_hd__and4_1_0/X CI sky130_fd_sc_hd__a21o_1_2/X
+ VNB VNB VPB VPB CO sky130_fd_sc_hd__a21o_1_3/a_384_47# sky130_fd_sc_hd__a21o_1_3/a_81_21#
+ sky130_fd_sc_hd__a21o_1_3/a_299_297# sky130_fd_sc_hd__a21o_1
Xsky130_fd_sc_hd__and4_1_0 P4 P2 P3 P1 VNB VNB VPB VPB sky130_fd_sc_hd__and4_1_0/X
+ sky130_fd_sc_hd__and4_1_0/a_109_47# sky130_fd_sc_hd__and4_1_0/a_197_47# sky130_fd_sc_hd__and4_1_0/a_303_47#
+ sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__and4_1
C0 CI VNB 0.02f
C1 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__a21o_1_0/X 0.00439f
C2 sky130_fd_sc_hd__a21o_1_2/X P2 0.455f
C3 sky130_fd_sc_hd__a21o_1_0/a_81_21# sky130_fd_sc_hd__a21o_1_2/X 8.44e-20
C4 G4 sky130_fd_sc_hd__a21o_1_1/X 0.0897f
C5 sky130_fd_sc_hd__and4_1_0/a_109_47# sky130_fd_sc_hd__and4_1_0/X 1.62e-19
C6 sky130_fd_sc_hd__a21o_1_1/a_299_297# P2 0.0566f
C7 G1 sky130_fd_sc_hd__a21o_1_1/X 0.00394f
C8 VNB sky130_fd_sc_hd__a21o_1_0/a_384_47# -2.71e-19
C9 sky130_fd_sc_hd__and4_1_0/a_109_47# VNB -6.28e-20
C10 P1 sky130_fd_sc_hd__a21o_1_1/X 4.83e-20
C11 sky130_fd_sc_hd__and4_1_0/a_27_47# VPB -0.0199f
C12 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__a21o_1_1/a_299_297# 0.0334f
C13 G1 sky130_fd_sc_hd__a21o_1_0/a_299_297# 0.0137f
C14 sky130_fd_sc_hd__and4_1_0/a_27_47# P3 0.0397f
C15 P3 VPB 0.0048f
C16 sky130_fd_sc_hd__and4_1_0/a_197_47# VPB -5.24e-19
C17 sky130_fd_sc_hd__a21o_1_1/a_384_47# VPB -4.08e-19
C18 sky130_fd_sc_hd__a21o_1_0/X sky130_fd_sc_hd__a21o_1_1/X 0.121f
C19 sky130_fd_sc_hd__and4_1_0/a_197_47# P3 0.0016f
C20 sky130_fd_sc_hd__and4_1_0/a_27_47# P4 0.00576f
C21 P2 sky130_fd_sc_hd__a21o_1_1/X 0.627f
C22 sky130_fd_sc_hd__a21o_1_0/a_81_21# sky130_fd_sc_hd__a21o_1_1/X 0.0018f
C23 G4 sky130_fd_sc_hd__and4_1_0/X 1.98e-20
C24 P3 sky130_fd_sc_hd__a21o_1_1/a_384_47# 7.45e-20
C25 sky130_fd_sc_hd__a21o_1_2/a_384_47# VPB -4.08e-19
C26 P4 VPB 0.0594f
C27 sky130_fd_sc_hd__a21o_1_2/a_81_21# VPB -0.0132f
C28 sky130_fd_sc_hd__a21o_1_2/a_384_47# P3 0.0013f
C29 P4 P3 0.2f
C30 P3 sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.0706f
C31 sky130_fd_sc_hd__a21o_1_0/X sky130_fd_sc_hd__a21o_1_0/a_299_297# 0.00259f
C32 G4 VNB 8.25e-19
C33 sky130_fd_sc_hd__a21o_1_1/a_81_21# VPB -0.00647f
C34 sky130_fd_sc_hd__a21o_1_0/a_299_297# P2 0.0456f
C35 CO P1 0.00943f
C36 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__a21o_1_1/X 0.0261f
C37 G3 VPB -6.71e-19
C38 P1 sky130_fd_sc_hd__and4_1_0/X 0.00732f
C39 sky130_fd_sc_hd__a21o_1_2/a_384_47# P4 6.19e-21
C40 P4 sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.00149f
C41 VNB G1 -0.00488f
C42 P3 G3 0.0176f
C43 sky130_fd_sc_hd__a21o_1_3/a_299_297# VPB -5.68e-32
C44 VPB sky130_fd_sc_hd__and4_1_0/a_303_47# -4.83e-19
C45 sky130_fd_sc_hd__a21o_1_1/a_299_297# sky130_fd_sc_hd__a21o_1_1/X 0.0338f
C46 VNB P1 0.0237f
C47 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__a21o_1_0/a_299_297# 1.65e-19
C48 P4 sky130_fd_sc_hd__a21o_1_1/a_81_21# 1.01e-19
C49 P3 sky130_fd_sc_hd__and4_1_0/a_303_47# 4.7e-19
C50 CO P2 4.84e-19
C51 sky130_fd_sc_hd__a21o_1_0/X sky130_fd_sc_hd__and4_1_0/X 7.95e-21
C52 sky130_fd_sc_hd__and4_1_0/X P2 0.00135f
C53 CI VPB 0.00996f
C54 sky130_fd_sc_hd__a21o_1_1/a_81_21# G3 0.023f
C55 VNB sky130_fd_sc_hd__a21o_1_0/X 0.461f
C56 VNB P2 0.00318f
C57 sky130_fd_sc_hd__a21o_1_0/a_81_21# VNB -0.0202f
C58 sky130_fd_sc_hd__a21o_1_2/X CO 0.0504f
C59 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__and4_1_0/X 0.132f
C60 P1 sky130_fd_sc_hd__a21o_1_3/a_81_21# 0.00196f
C61 sky130_fd_sc_hd__a21o_1_2/a_299_297# P2 0.055f
C62 sky130_fd_sc_hd__a21o_1_0/a_384_47# VPB -3.87e-19
C63 sky130_fd_sc_hd__and4_1_0/a_109_47# VPB -4.66e-19
C64 sky130_fd_sc_hd__a21o_1_2/X VNB 0.0224f
C65 G2 G1 0.0921f
C66 sky130_fd_sc_hd__and4_1_0/a_109_47# P3 0.00143f
C67 sky130_fd_sc_hd__a21o_1_0/a_299_297# sky130_fd_sc_hd__a21o_1_1/X 0.0315f
C68 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__a21o_1_2/a_299_297# 0.0335f
C69 CI sky130_fd_sc_hd__a21o_1_3/a_299_297# 0.00978f
C70 VNB sky130_fd_sc_hd__a21o_1_1/a_299_297# -0.00449f
C71 sky130_fd_sc_hd__a21o_1_3/a_81_21# P2 6.76e-19
C72 G2 sky130_fd_sc_hd__a21o_1_0/X 0.0575f
C73 G2 P2 0.00123f
C74 sky130_fd_sc_hd__a21o_1_0/a_81_21# G2 0.0401f
C75 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__a21o_1_3/a_81_21# 0.07f
C76 sky130_fd_sc_hd__and4_1_0/X sky130_fd_sc_hd__a21o_1_1/X 5.37e-20
C77 G4 VPB -0.00221f
C78 P3 G4 0.0694f
C79 VPB G1 0.0196f
C80 sky130_fd_sc_hd__a21o_1_2/X G2 5.09e-20
C81 VNB sky130_fd_sc_hd__a21o_1_1/X 0.0139f
C82 sky130_fd_sc_hd__and4_1_0/a_27_47# P1 0.019f
C83 G4 sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.0188f
C84 VPB P1 0.00652f
C85 P4 G4 0.02f
C86 sky130_fd_sc_hd__a21o_1_2/a_299_297# sky130_fd_sc_hd__a21o_1_1/X 0.0193f
C87 P3 P1 0.0581f
C88 VNB sky130_fd_sc_hd__a21o_1_0/a_299_297# -0.00449f
C89 sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__a21o_1_0/X 2.06e-20
C90 sky130_fd_sc_hd__and4_1_0/a_27_47# P2 0.0709f
C91 CO sky130_fd_sc_hd__and4_1_0/X 0.13f
C92 VPB sky130_fd_sc_hd__a21o_1_0/X 0.0377f
C93 sky130_fd_sc_hd__a21o_1_3/a_384_47# sky130_fd_sc_hd__and4_1_0/X 7.24e-19
C94 P4 P1 4.35e-19
C95 sky130_fd_sc_hd__a21o_1_2/a_81_21# P1 3.15e-20
C96 VPB P2 0.383f
C97 sky130_fd_sc_hd__a21o_1_0/a_81_21# VPB -0.00151f
C98 P3 sky130_fd_sc_hd__a21o_1_0/X 0.0694f
C99 sky130_fd_sc_hd__and4_1_0/a_197_47# sky130_fd_sc_hd__a21o_1_0/X 5.93e-21
C100 P3 P2 0.155f
C101 sky130_fd_sc_hd__and4_1_0/a_197_47# P2 2.63e-19
C102 sky130_fd_sc_hd__a21o_1_1/a_384_47# sky130_fd_sc_hd__a21o_1_0/X 6.97e-19
C103 VNB sky130_fd_sc_hd__a21o_1_3/a_384_47# -5.85e-20
C104 CO VNB -0.00689f
C105 VNB sky130_fd_sc_hd__and4_1_0/X 0.251f
C106 sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__a21o_1_2/X 0.0588f
C107 G3 P1 3.23e-21
C108 sky130_fd_sc_hd__a21o_1_2/a_384_47# sky130_fd_sc_hd__a21o_1_0/X 1.12e-20
C109 sky130_fd_sc_hd__a21o_1_2/a_81_21# sky130_fd_sc_hd__a21o_1_0/X 1.2e-19
C110 P4 sky130_fd_sc_hd__a21o_1_0/X 5.9e-20
C111 sky130_fd_sc_hd__a21o_1_2/X VPB 1.21f
C112 sky130_fd_sc_hd__a21o_1_2/a_384_47# P2 2.47e-20
C113 P4 P2 0.197f
C114 sky130_fd_sc_hd__a21o_1_2/a_81_21# P2 0.0301f
C115 G2 sky130_fd_sc_hd__a21o_1_1/X 1.59e-19
C116 sky130_fd_sc_hd__a21o_1_3/a_299_297# P1 2.61e-19
C117 P3 sky130_fd_sc_hd__a21o_1_2/X 0.0674f
C118 sky130_fd_sc_hd__a21o_1_1/a_81_21# sky130_fd_sc_hd__a21o_1_0/X 0.0631f
C119 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__a21o_1_1/a_384_47# 1.32e-20
C120 sky130_fd_sc_hd__a21o_1_1/a_81_21# P2 0.0526f
C121 G3 sky130_fd_sc_hd__a21o_1_0/X 0.0894f
C122 VPB sky130_fd_sc_hd__a21o_1_1/a_299_297# -0.00193f
C123 G3 P2 0.0287f
C124 CI P1 2.89e-19
C125 P4 sky130_fd_sc_hd__a21o_1_2/X 0.00977f
C126 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.02f
C127 VNB sky130_fd_sc_hd__a21o_1_2/a_299_297# -0.00449f
C128 P3 sky130_fd_sc_hd__a21o_1_1/a_299_297# 0.00415f
C129 CO sky130_fd_sc_hd__a21o_1_3/a_81_21# 0.00936f
C130 sky130_fd_sc_hd__a21o_1_0/X sky130_fd_sc_hd__and4_1_0/a_303_47# 5.18e-21
C131 sky130_fd_sc_hd__and4_1_0/X sky130_fd_sc_hd__a21o_1_3/a_81_21# 0.0697f
C132 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__a21o_1_1/a_81_21# 0.00223f
C133 P4 sky130_fd_sc_hd__a21o_1_1/a_299_297# 1.23e-19
C134 sky130_fd_sc_hd__a21o_1_2/X G3 4.15e-19
C135 sky130_fd_sc_hd__a21o_1_0/a_384_47# G1 4.61e-19
C136 VNB sky130_fd_sc_hd__a21o_1_3/a_81_21# -0.0199f
C137 CI P2 2.97e-20
C138 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__a21o_1_3/a_299_297# 0.0173f
C139 sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__a21o_1_1/X 1.67e-19
C140 sky130_fd_sc_hd__a21o_1_2/X sky130_fd_sc_hd__and4_1_0/a_303_47# 4.26e-19
C141 VPB sky130_fd_sc_hd__a21o_1_1/X 0.0255f
C142 P3 sky130_fd_sc_hd__a21o_1_1/X 0.185f
C143 VNB G2 0.00126f
C144 sky130_fd_sc_hd__a21o_1_2/X CI 0.00156f
C145 sky130_fd_sc_hd__a21o_1_1/a_384_47# sky130_fd_sc_hd__a21o_1_1/X 4.81e-19
C146 sky130_fd_sc_hd__a21o_1_0/a_384_47# sky130_fd_sc_hd__a21o_1_0/X 0.00135f
C147 sky130_fd_sc_hd__and4_1_0/a_109_47# sky130_fd_sc_hd__a21o_1_0/X 9.17e-21
C148 VPB sky130_fd_sc_hd__a21o_1_0/a_299_297# 0.00347f
C149 sky130_fd_sc_hd__and4_1_0/a_109_47# P2 2.77e-19
C150 sky130_fd_sc_hd__a21o_1_2/a_384_47# sky130_fd_sc_hd__a21o_1_1/X 7.94e-20
C151 P4 sky130_fd_sc_hd__a21o_1_1/X 0.0428f
C152 sky130_fd_sc_hd__a21o_1_2/a_81_21# sky130_fd_sc_hd__a21o_1_1/X 0.0421f
C153 sky130_fd_sc_hd__a21o_1_1/a_81_21# sky130_fd_sc_hd__a21o_1_1/X 0.0447f
C154 sky130_fd_sc_hd__and4_1_0/a_27_47# CO 0.00246f
C155 G3 sky130_fd_sc_hd__a21o_1_1/X 0.0595f
C156 G4 P1 1.7e-20
C157 sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__and4_1_0/X 0.00169f
C158 CO VPB -0.00363f
C159 VPB sky130_fd_sc_hd__a21o_1_3/a_384_47# -1.62e-19
C160 VPB sky130_fd_sc_hd__and4_1_0/X 0.0202f
C161 P3 CO 0.0012f
C162 P3 sky130_fd_sc_hd__and4_1_0/X 0.00586f
C163 sky130_fd_sc_hd__and4_1_0/a_197_47# sky130_fd_sc_hd__and4_1_0/X 1.78e-19
C164 sky130_fd_sc_hd__and4_1_0/a_27_47# VNB 0.00805f
C165 sky130_fd_sc_hd__a21o_1_1/a_384_47# sky130_fd_sc_hd__and4_1_0/X 1.46e-21
C166 VNB VPB -0.275f
C167 G4 sky130_fd_sc_hd__a21o_1_0/X 3.47e-20
C168 G4 P2 0.00574f
C169 sky130_fd_sc_hd__a21o_1_2/a_384_47# sky130_fd_sc_hd__and4_1_0/X 1.23e-20
C170 P4 sky130_fd_sc_hd__and4_1_0/X 4.68e-20
C171 sky130_fd_sc_hd__a21o_1_2/a_81_21# sky130_fd_sc_hd__and4_1_0/X 4.69e-20
C172 P3 VNB 0.543f
C173 sky130_fd_sc_hd__and4_1_0/a_197_47# VNB -4.52e-20
C174 sky130_fd_sc_hd__a21o_1_1/a_384_47# VNB -1.89e-19
C175 G1 sky130_fd_sc_hd__a21o_1_0/X 0.0691f
C176 VPB sky130_fd_sc_hd__a21o_1_2/a_299_297# 0.0196f
C177 G1 P2 0.0935f
C178 sky130_fd_sc_hd__a21o_1_0/a_81_21# G1 0.00416f
C179 sky130_fd_sc_hd__a21o_1_2/a_384_47# VNB -2.27e-19
C180 P3 sky130_fd_sc_hd__a21o_1_2/a_299_297# 0.00159f
C181 P4 VNB 0.00496f
C182 sky130_fd_sc_hd__a21o_1_2/a_81_21# VNB -0.0181f
C183 P1 sky130_fd_sc_hd__a21o_1_0/X 1.23e-20
C184 sky130_fd_sc_hd__a21o_1_2/X G4 0.00776f
C185 P1 P2 0.0215f
C186 sky130_fd_sc_hd__and4_1_0/a_27_47# sky130_fd_sc_hd__a21o_1_3/a_81_21# 0.0108f
C187 sky130_fd_sc_hd__a21o_1_0/a_384_47# sky130_fd_sc_hd__a21o_1_1/X 1.32e-20
C188 sky130_fd_sc_hd__a21o_1_3/a_299_297# sky130_fd_sc_hd__and4_1_0/X 0.00642f
C189 sky130_fd_sc_hd__a21o_1_1/a_81_21# VNB -0.0191f
C190 P4 sky130_fd_sc_hd__a21o_1_2/a_299_297# 0.0108f
C191 sky130_fd_sc_hd__a21o_1_2/X G1 4.98e-20
C192 VPB sky130_fd_sc_hd__a21o_1_3/a_81_21# -0.0123f
C193 sky130_fd_sc_hd__and4_1_0/X sky130_fd_sc_hd__and4_1_0/a_303_47# 3.17e-19
C194 G3 VNB 6.81e-19
C195 P3 sky130_fd_sc_hd__a21o_1_3/a_81_21# 2.3e-19
C196 sky130_fd_sc_hd__a21o_1_2/X P1 0.0247f
C197 sky130_fd_sc_hd__a21o_1_0/X P2 0.0752f
C198 sky130_fd_sc_hd__a21o_1_0/a_81_21# sky130_fd_sc_hd__a21o_1_0/X 0.059f
C199 sky130_fd_sc_hd__a21o_1_3/a_299_297# VNB -0.00378f
C200 sky130_fd_sc_hd__a21o_1_0/a_81_21# P2 0.00281f
C201 CI sky130_fd_sc_hd__and4_1_0/X 0.0308f
C202 VNB sky130_fd_sc_hd__and4_1_0/a_303_47# 3.12e-20
C203 VPB G2 0.0175f
C204 VNB 0 1.71f
C205 VPB 0 4.61f
C206 sky130_fd_sc_hd__and4_1_0/X 0 0.154f
C207 P1 0 0.164f
C208 P3 0 0.297f
C209 P2 0 0.31f
C210 P4 0 0.324f
C211 sky130_fd_sc_hd__and4_1_0/a_27_47# 0 0.175f
C212 CO 0 0.0276f
C213 CI 0 0.158f
C214 sky130_fd_sc_hd__a21o_1_3/a_299_297# 0 0.0348f
C215 sky130_fd_sc_hd__a21o_1_3/a_81_21# 0 0.147f
C216 sky130_fd_sc_hd__a21o_1_2/X 0 0.168f
C217 sky130_fd_sc_hd__a21o_1_1/X 0 0.129f
C218 G4 0 0.137f
C219 sky130_fd_sc_hd__a21o_1_2/a_299_297# 0 0.0348f
C220 sky130_fd_sc_hd__a21o_1_2/a_81_21# 0 0.147f
C221 sky130_fd_sc_hd__a21o_1_0/X 0 0.223f
C222 G3 0 0.137f
C223 sky130_fd_sc_hd__a21o_1_1/a_299_297# 0 0.0348f
C224 sky130_fd_sc_hd__a21o_1_1/a_81_21# 0 0.147f
C225 G1 0 0.12f
C226 G2 0 0.163f
C227 sky130_fd_sc_hd__a21o_1_0/a_299_297# 0 0.0348f
C228 sky130_fd_sc_hd__a21o_1_0/a_81_21# 0 0.147f
.ends

.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X a_117_297# a_285_297# a_285_47#
+ a_35_297#
X0 X a_35_297# a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.177 ps=1.69 w=1 l=0.15
**devattr s=10400,504 d=12000,520
X1 X B a_285_47# VNB sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.42 as=0.0878 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=10010,284
X2 a_35_297# B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.138 ps=1.4 w=0.65 l=0.15
**devattr s=6760,364 d=3510,184
X3 a_117_297# B a_35_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
**devattr s=10400,504 d=5400,254
X4 VPWR B a_285_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.177 pd=1.69 as=0.177 ps=1.69 w=1 l=0.15
**devattr s=5400,254 d=10400,504
X5 VGND A a_35_297# VNB sky130_fd_pr__nfet_01v8 ad=0.138 pd=1.4 as=0.0878 ps=0.92 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
X6 VGND a_35_297# X VNB sky130_fd_pr__nfet_01v8 ad=0.138 pd=1.4 as=0.25 ps=1.42 w=0.65 l=0.15
**devattr s=10010,284 d=8320,388
X7 a_285_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.177 pd=1.69 as=0.177 ps=1.69 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X8 VPWR A a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.177 pd=1.69 as=0.135 ps=1.27 w=1 l=0.15
**devattr s=5400,254 d=5400,254
X9 a_285_47# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.92 as=0.138 ps=1.4 w=0.65 l=0.15
**devattr s=3510,184 d=3510,184
C0 a_285_297# VPB 0.0133f
C1 a_117_297# X 2.25e-19
C2 VGND VPB 0.00696f
C3 B VPB 0.0697f
C4 a_35_297# A 0.0633f
C5 a_35_297# a_285_297# 0.025f
C6 a_35_297# VGND 0.177f
C7 a_35_297# B 0.203f
C8 a_35_297# VPB 0.0699f
C9 a_285_47# VGND 0.00552f
C10 X VPWR 0.0537f
C11 a_285_47# B 3.98e-19
C12 a_117_297# VGND 0.00177f
C13 a_117_297# B 0.00777f
C14 a_35_297# a_285_47# 0.00723f
C15 A VPWR 0.0348f
C16 a_285_297# VPWR 0.246f
C17 a_117_297# a_35_297# 0.00641f
C18 VGND VPWR 0.0643f
C19 B VPWR 0.0703f
C20 A X 0.00166f
C21 a_285_297# X 0.0712f
C22 VPWR VPB 0.0689f
C23 X VGND 0.173f
C24 X B 0.0149f
C25 a_35_297# VPWR 0.096f
C26 X VPB 0.0154f
C27 a_285_47# VPWR 8.6e-19
C28 a_35_297# X 0.166f
C29 a_285_297# A 0.00749f
C30 A VGND 0.0325f
C31 A B 0.221f
C32 a_285_297# VGND 0.00394f
C33 a_285_297# B 0.0553f
C34 a_117_297# VPWR 0.00852f
C35 X a_285_47# 0.00206f
C36 VGND B 0.0304f
C37 A VPB 0.051f
C38 VGND VNB 0.435f
C39 X VNB 0.0649f
C40 VPWR VNB 0.333f
C41 A VNB 0.167f
C42 B VNB 0.213f
C43 VPB VNB 0.693f
C44 a_285_297# VNB 0.00137f
C45 a_35_297# VNB 0.255f
.ends

.subckt adder_3 G1 P2 G2 G3 P4 S1 S2 S3 S4 sky130_fd_sc_hd__xor2_1_3/a_117_297# sky130_fd_sc_hd__xor2_1_3/a_35_297#
+ sky130_fd_sc_hd__a21o_1_0/a_81_21# sky130_fd_sc_hd__xor2_1_3/a_285_47# sky130_fd_sc_hd__xor2_1_0/a_285_297#
+ sky130_fd_sc_hd__a21o_1_0/a_384_47# sky130_fd_sc_hd__xor2_1_1/a_285_297# sky130_fd_sc_hd__xor2_1_0/a_35_297#
+ sky130_fd_sc_hd__xor2_1_0/a_285_47# sky130_fd_sc_hd__a21o_1_1/a_81_21# sky130_fd_sc_hd__a21o_1_0/a_299_297#
+ sky130_fd_sc_hd__xor2_1_2/a_285_297# sky130_fd_sc_hd__xor2_1_3/a_285_297# sky130_fd_sc_hd__a21o_1_1/a_299_297#
+ sky130_fd_sc_hd__a21o_1_2/a_299_297# sky130_fd_sc_hd__xor2_1_1/a_35_297# sky130_fd_sc_hd__xor2_1_3/B
+ sky130_fd_sc_hd__xor2_1_1/a_285_47# sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__a21o_1_2/a_81_21#
+ sky130_fd_sc_hd__xor2_1_0/a_117_297# sky130_fd_sc_hd__xor2_1_2/a_35_297# sky130_fd_sc_hd__xor2_1_2/a_285_47#
+ sky130_fd_sc_hd__xor2_1_1/a_117_297# CI P1 SUB sky130_fd_sc_hd__xor2_1_2/B sky130_fd_sc_hd__xor2_1_2/a_117_297#
+ VPB P3
Xsky130_fd_sc_hd__xor2_1_3 P4 sky130_fd_sc_hd__xor2_1_3/B SUB SUB VPB VPB S4 sky130_fd_sc_hd__xor2_1_3/a_117_297#
+ sky130_fd_sc_hd__xor2_1_3/a_285_297# sky130_fd_sc_hd__xor2_1_3/a_285_47# sky130_fd_sc_hd__xor2_1_3/a_35_297#
+ sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__a21o_1_0 CI P1 G1 SUB SUB VPB VPB sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__a21o_1_0/a_384_47#
+ sky130_fd_sc_hd__a21o_1_0/a_81_21# sky130_fd_sc_hd__a21o_1_0/a_299_297# sky130_fd_sc_hd__a21o_1
Xsky130_fd_sc_hd__a21o_1_1 sky130_fd_sc_hd__xor2_1_1/B P2 G2 SUB SUB VPB VPB sky130_fd_sc_hd__xor2_1_2/B
+ sky130_fd_sc_hd__a21o_1_1/a_384_47# sky130_fd_sc_hd__a21o_1_1/a_81_21# sky130_fd_sc_hd__a21o_1_1/a_299_297#
+ sky130_fd_sc_hd__a21o_1
Xsky130_fd_sc_hd__a21o_1_2 sky130_fd_sc_hd__xor2_1_2/B P3 G3 SUB SUB VPB VPB sky130_fd_sc_hd__xor2_1_3/B
+ sky130_fd_sc_hd__a21o_1_2/a_384_47# sky130_fd_sc_hd__a21o_1_2/a_81_21# sky130_fd_sc_hd__a21o_1_2/a_299_297#
+ sky130_fd_sc_hd__a21o_1
Xsky130_fd_sc_hd__xor2_1_0 P1 CI SUB SUB VPB VPB S1 sky130_fd_sc_hd__xor2_1_0/a_117_297#
+ sky130_fd_sc_hd__xor2_1_0/a_285_297# sky130_fd_sc_hd__xor2_1_0/a_285_47# sky130_fd_sc_hd__xor2_1_0/a_35_297#
+ sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_1 P2 sky130_fd_sc_hd__xor2_1_1/B SUB SUB VPB VPB S2 sky130_fd_sc_hd__xor2_1_1/a_117_297#
+ sky130_fd_sc_hd__xor2_1_1/a_285_297# sky130_fd_sc_hd__xor2_1_1/a_285_47# sky130_fd_sc_hd__xor2_1_1/a_35_297#
+ sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_2 P3 sky130_fd_sc_hd__xor2_1_2/B SUB SUB VPB VPB S3 sky130_fd_sc_hd__xor2_1_2/a_117_297#
+ sky130_fd_sc_hd__xor2_1_2/a_285_297# sky130_fd_sc_hd__xor2_1_2/a_285_47# sky130_fd_sc_hd__xor2_1_2/a_35_297#
+ sky130_fd_sc_hd__xor2_1
C0 P2 G3 0.0223f
C1 VPB sky130_fd_sc_hd__xor2_1_2/a_285_297# 2.35e-20
C2 S3 sky130_fd_sc_hd__xor2_1_2/a_117_297# 6.67e-19
C3 sky130_fd_sc_hd__xor2_1_1/a_35_297# sky130_fd_sc_hd__xor2_1_2/B 0.0151f
C4 S3 sky130_fd_sc_hd__xor2_1_3/a_35_297# 0.0518f
C5 sky130_fd_sc_hd__a21o_1_2/a_299_297# S1 3.56e-19
C6 P2 SUB 0.384f
C7 sky130_fd_sc_hd__xor2_1_0/a_285_47# P1 0.00118f
C8 sky130_fd_sc_hd__a21o_1_2/a_384_47# sky130_fd_sc_hd__xor2_1_2/B 0.00105f
C9 S2 sky130_fd_sc_hd__xor2_1_1/a_285_297# 0.00293f
C10 sky130_fd_sc_hd__xor2_1_3/a_285_47# sky130_fd_sc_hd__xor2_1_3/B 3.65e-19
C11 S3 sky130_fd_sc_hd__xor2_1_1/a_35_297# 3.35e-20
C12 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__a21o_1_0/a_384_47# 3.85e-19
C13 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__a21o_1_1/a_384_47# 0.00123f
C14 G3 sky130_fd_sc_hd__xor2_1_3/B 0.0517f
C15 sky130_fd_sc_hd__xor2_1_1/a_35_297# P1 0.00101f
C16 sky130_fd_sc_hd__xor2_1_1/B VPB 0.743f
C17 P3 S1 2.04e-19
C18 sky130_fd_sc_hd__xor2_1_3/B SUB 1.3f
C19 CI S1 0.002f
C20 P2 sky130_fd_sc_hd__xor2_1_3/B 0.107f
C21 sky130_fd_sc_hd__a21o_1_2/a_81_21# S1 2.24e-19
C22 VPB sky130_fd_sc_hd__xor2_1_0/a_117_297# -2.04e-19
C23 P4 P3 4.73e-19
C24 sky130_fd_sc_hd__xor2_1_2/a_35_297# S2 0.0515f
C25 sky130_fd_sc_hd__xor2_1_3/a_117_297# S4 6.67e-19
C26 G3 sky130_fd_sc_hd__xor2_1_2/B 0.0811f
C27 sky130_fd_sc_hd__xor2_1_2/a_285_297# S2 0.00111f
C28 sky130_fd_sc_hd__a21o_1_1/a_299_297# S1 8.32e-20
C29 SUB sky130_fd_sc_hd__xor2_1_2/B 0.233f
C30 P2 sky130_fd_sc_hd__xor2_1_2/B 0.163f
C31 sky130_fd_sc_hd__xor2_1_1/B G2 0.13f
C32 G3 P1 6.62e-19
C33 S3 SUB -0.00162f
C34 sky130_fd_sc_hd__a21o_1_0/a_299_297# SUB -0.00435f
C35 S3 P2 2.48e-20
C36 sky130_fd_sc_hd__xor2_1_0/a_35_297# P3 0.00793f
C37 sky130_fd_sc_hd__xor2_1_1/B S2 0.00554f
C38 P1 SUB 1f
C39 sky130_fd_sc_hd__xor2_1_3/a_35_297# sky130_fd_sc_hd__xor2_1_2/a_35_297# 0.00123f
C40 CI sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.0235f
C41 sky130_fd_sc_hd__xor2_1_3/B sky130_fd_sc_hd__xor2_1_2/B 0.171f
C42 sky130_fd_sc_hd__a21o_1_2/a_81_21# sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.00109f
C43 P2 P1 0.6f
C44 VPB sky130_fd_sc_hd__a21o_1_2/a_299_297# 0.0344f
C45 sky130_fd_sc_hd__xor2_1_1/a_35_297# sky130_fd_sc_hd__xor2_1_2/a_35_297# 0.00123f
C46 S3 sky130_fd_sc_hd__xor2_1_3/B 0.0617f
C47 VPB sky130_fd_sc_hd__xor2_1_2/a_285_47# -7.24e-19
C48 CI sky130_fd_sc_hd__a21o_1_0/a_384_47# 0.00162f
C49 sky130_fd_sc_hd__xor2_1_3/B P1 0.0733f
C50 VPB P3 0.0315f
C51 P4 S4 0.00239f
C52 sky130_fd_sc_hd__xor2_1_3/a_285_297# S4 0.00453f
C53 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__xor2_1_0/a_285_47# 2.47e-19
C54 VPB CI 0.00219f
C55 VPB sky130_fd_sc_hd__a21o_1_2/a_81_21# -0.00306f
C56 SUB sky130_fd_sc_hd__xor2_1_1/a_285_297# -0.00394f
C57 S3 sky130_fd_sc_hd__xor2_1_2/B 0.00532f
C58 sky130_fd_sc_hd__a21o_1_0/a_299_297# sky130_fd_sc_hd__xor2_1_2/B 0.0414f
C59 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__xor2_1_3/a_35_297# 5.05e-21
C60 VPB sky130_fd_sc_hd__a21o_1_0/a_81_21# -0.00793f
C61 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.0394f
C62 P1 sky130_fd_sc_hd__xor2_1_2/B 0.183f
C63 VPB sky130_fd_sc_hd__a21o_1_1/a_299_297# 0.0016f
C64 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__a21o_1_2/a_384_47# 2.81e-20
C65 sky130_fd_sc_hd__a21o_1_0/a_299_297# P1 0.00669f
C66 sky130_fd_sc_hd__xor2_1_3/B sky130_fd_sc_hd__xor2_1_1/a_285_297# 0.00704f
C67 sky130_fd_sc_hd__xor2_1_2/a_35_297# SUB -0.0113f
C68 P2 sky130_fd_sc_hd__xor2_1_2/a_35_297# 6.69e-19
C69 CI G2 2.73e-19
C70 sky130_fd_sc_hd__xor2_1_2/a_285_297# SUB -0.00394f
C71 S2 P3 0.00112f
C72 sky130_fd_sc_hd__a21o_1_0/a_81_21# G2 1.77e-20
C73 VPB sky130_fd_sc_hd__a21o_1_1/a_81_21# -0.00424f
C74 sky130_fd_sc_hd__xor2_1_1/B G3 0.0538f
C75 sky130_fd_sc_hd__xor2_1_3/B sky130_fd_sc_hd__xor2_1_2/a_35_297# 0.0908f
C76 VPB G1 0.00163f
C77 S3 sky130_fd_sc_hd__xor2_1_1/a_285_297# 8.64e-20
C78 VPB S4 0.0296f
C79 sky130_fd_sc_hd__xor2_1_2/a_285_297# sky130_fd_sc_hd__xor2_1_3/B 0.00704f
C80 sky130_fd_sc_hd__xor2_1_1/B SUB 0.137f
C81 sky130_fd_sc_hd__xor2_1_1/B P2 0.223f
C82 sky130_fd_sc_hd__xor2_1_2/a_35_297# sky130_fd_sc_hd__xor2_1_2/B 0.0262f
C83 SUB sky130_fd_sc_hd__xor2_1_0/a_117_297# -0.00177f
C84 sky130_fd_sc_hd__xor2_1_3/a_35_297# P3 0.00203f
C85 G2 sky130_fd_sc_hd__a21o_1_1/a_81_21# 0.0275f
C86 S3 sky130_fd_sc_hd__xor2_1_2/a_35_297# 0.00495f
C87 sky130_fd_sc_hd__xor2_1_1/a_35_297# P3 2.02e-19
C88 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__xor2_1_3/B 0.398f
C89 G1 G2 1.42e-20
C90 CI sky130_fd_sc_hd__xor2_1_1/a_35_297# 7.26e-21
C91 S3 sky130_fd_sc_hd__xor2_1_2/a_285_297# 0.00453f
C92 sky130_fd_sc_hd__a21o_1_2/a_384_47# P3 5.7e-19
C93 VPB sky130_fd_sc_hd__xor2_1_3/a_117_297# 2.25e-20
C94 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__xor2_1_2/B 0.161f
C95 VPB sky130_fd_sc_hd__xor2_1_1/a_285_47# -7.24e-19
C96 sky130_fd_sc_hd__xor2_1_3/a_285_47# P3 3.53e-19
C97 sky130_fd_sc_hd__xor2_1_0/a_285_297# S1 0.00385f
C98 sky130_fd_sc_hd__xor2_1_1/B S3 3.34e-20
C99 sky130_fd_sc_hd__xor2_1_0/a_117_297# sky130_fd_sc_hd__xor2_1_2/B 2.27e-19
C100 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__a21o_1_0/a_299_297# 0.0526f
C101 sky130_fd_sc_hd__a21o_1_2/a_299_297# SUB -0.00449f
C102 sky130_fd_sc_hd__xor2_1_0/a_35_297# S1 0.00396f
C103 sky130_fd_sc_hd__xor2_1_1/a_117_297# S1 0.00102f
C104 sky130_fd_sc_hd__xor2_1_2/a_285_47# SUB -4.65e-19
C105 sky130_fd_sc_hd__xor2_1_1/B P1 0.132f
C106 CI G3 2.35e-19
C107 G3 sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.0232f
C108 SUB P3 0.27f
C109 P2 P3 0.608f
C110 sky130_fd_sc_hd__a21o_1_2/a_299_297# sky130_fd_sc_hd__xor2_1_3/B 6.06e-19
C111 CI SUB 0.176f
C112 sky130_fd_sc_hd__xor2_1_3/a_35_297# S4 0.00521f
C113 sky130_fd_sc_hd__a21o_1_2/a_81_21# SUB -0.0181f
C114 CI P2 0.186f
C115 P2 sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.0197f
C116 sky130_fd_sc_hd__xor2_1_2/a_285_47# sky130_fd_sc_hd__xor2_1_3/B 0.00259f
C117 sky130_fd_sc_hd__a21o_1_0/a_81_21# SUB -0.00347f
C118 VPB S1 0.0368f
C119 sky130_fd_sc_hd__a21o_1_1/a_299_297# SUB -0.00436f
C120 sky130_fd_sc_hd__xor2_1_3/B P3 0.159f
C121 P2 sky130_fd_sc_hd__a21o_1_1/a_299_297# 0.00664f
C122 sky130_fd_sc_hd__a21o_1_2/a_299_297# sky130_fd_sc_hd__xor2_1_2/B 0.00554f
C123 CI sky130_fd_sc_hd__xor2_1_3/B 0.0784f
C124 VPB P4 0.0224f
C125 sky130_fd_sc_hd__xor2_1_3/B sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.0563f
C126 sky130_fd_sc_hd__a21o_1_0/a_81_21# sky130_fd_sc_hd__xor2_1_3/B 1.96e-19
C127 P3 sky130_fd_sc_hd__xor2_1_2/B 0.902f
C128 sky130_fd_sc_hd__xor2_1_3/B sky130_fd_sc_hd__a21o_1_1/a_299_297# 0.0322f
C129 CI sky130_fd_sc_hd__xor2_1_2/B 0.818f
C130 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__xor2_1_2/a_35_297# 6.93e-20
C131 sky130_fd_sc_hd__a21o_1_2/a_81_21# sky130_fd_sc_hd__xor2_1_2/B 0.0116f
C132 VPB sky130_fd_sc_hd__xor2_1_0/a_285_297# -3.91e-19
C133 SUB sky130_fd_sc_hd__a21o_1_1/a_81_21# -0.00243f
C134 S3 P3 0.00706f
C135 P2 sky130_fd_sc_hd__a21o_1_1/a_81_21# 0.00611f
C136 G1 SUB 0.023f
C137 VPB sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.042f
C138 sky130_fd_sc_hd__a21o_1_0/a_81_21# sky130_fd_sc_hd__xor2_1_2/B 0.00447f
C139 VPB sky130_fd_sc_hd__xor2_1_1/a_117_297# 2.29e-20
C140 sky130_fd_sc_hd__a21o_1_0/a_299_297# CI 0.00517f
C141 SUB S4 0.0195f
C142 sky130_fd_sc_hd__a21o_1_1/a_299_297# sky130_fd_sc_hd__xor2_1_2/B 0.00516f
C143 P1 P3 0.0282f
C144 S2 S1 0.0103f
C145 CI P1 0.544f
C146 sky130_fd_sc_hd__a21o_1_2/a_81_21# P1 2.85e-19
C147 sky130_fd_sc_hd__xor2_1_3/B sky130_fd_sc_hd__a21o_1_1/a_81_21# 0.00303f
C148 VPB sky130_fd_sc_hd__a21o_1_0/a_384_47# -4.08e-19
C149 G1 sky130_fd_sc_hd__xor2_1_3/B 1.88e-20
C150 sky130_fd_sc_hd__a21o_1_0/a_81_21# P1 7.84e-20
C151 VPB sky130_fd_sc_hd__a21o_1_1/a_384_47# -4.08e-19
C152 sky130_fd_sc_hd__xor2_1_3/B S4 0.00601f
C153 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__xor2_1_0/a_117_297# 0.00427f
C154 sky130_fd_sc_hd__xor2_1_2/a_117_297# S1 2.46e-20
C155 sky130_fd_sc_hd__a21o_1_1/a_81_21# sky130_fd_sc_hd__xor2_1_2/B 0.0211f
C156 G1 sky130_fd_sc_hd__xor2_1_2/B 0.0014f
C157 sky130_fd_sc_hd__xor2_1_3/a_117_297# SUB -8.18e-19
C158 sky130_fd_sc_hd__xor2_1_1/a_117_297# S2 5.82e-19
C159 sky130_fd_sc_hd__xor2_1_1/a_35_297# S1 0.0535f
C160 sky130_fd_sc_hd__xor2_1_3/a_35_297# P4 0.0132f
C161 sky130_fd_sc_hd__xor2_1_1/a_285_47# SUB -4.65e-19
C162 P2 sky130_fd_sc_hd__xor2_1_1/a_285_47# 0.00118f
C163 S3 S4 0.0102f
C164 P1 sky130_fd_sc_hd__a21o_1_1/a_81_21# 0.0152f
C165 sky130_fd_sc_hd__xor2_1_2/a_35_297# P3 0.0152f
C166 VPB G2 0.00129f
C167 sky130_fd_sc_hd__xor2_1_3/B sky130_fd_sc_hd__xor2_1_3/a_117_297# 0.00267f
C168 VPB S2 0.0397f
C169 sky130_fd_sc_hd__xor2_1_3/B sky130_fd_sc_hd__xor2_1_1/a_285_47# 0.00253f
C170 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__a21o_1_2/a_299_297# 0.0519f
C171 G3 S1 8.29e-20
C172 sky130_fd_sc_hd__xor2_1_1/a_35_297# sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.00128f
C173 sky130_fd_sc_hd__xor2_1_1/B P3 0.051f
C174 sky130_fd_sc_hd__xor2_1_1/a_285_47# sky130_fd_sc_hd__xor2_1_2/B 5.8e-19
C175 SUB S1 -0.00328f
C176 sky130_fd_sc_hd__a21o_1_2/a_384_47# sky130_fd_sc_hd__xor2_1_0/a_35_297# 6.06e-21
C177 S3 sky130_fd_sc_hd__xor2_1_3/a_117_297# 0.00101f
C178 P2 S1 0.00354f
C179 sky130_fd_sc_hd__xor2_1_1/B CI 0.155f
C180 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.0491f
C181 VPB sky130_fd_sc_hd__xor2_1_2/a_117_297# 2.25e-20
C182 VPB sky130_fd_sc_hd__xor2_1_0/a_285_47# -8.6e-19
C183 P4 SUB 0.0233f
C184 VPB sky130_fd_sc_hd__xor2_1_3/a_35_297# 0.00512f
C185 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__a21o_1_0/a_81_21# 0.0562f
C186 CI sky130_fd_sc_hd__xor2_1_0/a_117_297# 9.44e-19
C187 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__a21o_1_1/a_299_297# 0.0587f
C188 VPB sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.00693f
C189 sky130_fd_sc_hd__xor2_1_3/B S1 0.0317f
C190 G3 sky130_fd_sc_hd__xor2_1_0/a_35_297# 6.72e-20
C191 VPB sky130_fd_sc_hd__a21o_1_2/a_384_47# -4.08e-19
C192 SUB sky130_fd_sc_hd__xor2_1_0/a_285_297# -0.00394f
C193 P4 sky130_fd_sc_hd__xor2_1_3/B 0.104f
C194 SUB sky130_fd_sc_hd__xor2_1_0/a_35_297# -0.0143f
C195 sky130_fd_sc_hd__xor2_1_1/a_117_297# SUB -0.00177f
C196 sky130_fd_sc_hd__xor2_1_2/B S1 1.38e-19
C197 P2 sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.00129f
C198 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__a21o_1_1/a_81_21# 0.0601f
C199 sky130_fd_sc_hd__a21o_1_2/a_299_297# P3 0.00623f
C200 S3 S1 3.29e-19
C201 sky130_fd_sc_hd__xor2_1_2/a_117_297# S2 8.82e-19
C202 sky130_fd_sc_hd__xor2_1_1/B G1 0.0614f
C203 sky130_fd_sc_hd__xor2_1_3/B sky130_fd_sc_hd__xor2_1_0/a_285_297# 1.77e-19
C204 VPB G3 0.00152f
C205 sky130_fd_sc_hd__xor2_1_2/a_285_47# P3 0.00118f
C206 sky130_fd_sc_hd__a21o_1_0/a_384_47# SUB 4.44e-34
C207 sky130_fd_sc_hd__xor2_1_3/B sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.0707f
C208 sky130_fd_sc_hd__xor2_1_1/a_117_297# sky130_fd_sc_hd__xor2_1_3/B 0.00134f
C209 S3 P4 0.00111f
C210 P1 S1 0.00593f
C211 S3 sky130_fd_sc_hd__xor2_1_3/a_285_297# 0.00135f
C212 P2 sky130_fd_sc_hd__a21o_1_1/a_384_47# 6.47e-19
C213 sky130_fd_sc_hd__xor2_1_1/a_35_297# S2 0.00476f
C214 VPB SUB -0.376f
C215 VPB P2 0.0257f
C216 CI P3 0.346f
C217 sky130_fd_sc_hd__a21o_1_2/a_81_21# P3 4.57e-20
C218 CI sky130_fd_sc_hd__a21o_1_2/a_81_21# 1.2e-19
C219 sky130_fd_sc_hd__xor2_1_0/a_35_297# sky130_fd_sc_hd__xor2_1_2/B 0.00271f
C220 sky130_fd_sc_hd__xor2_1_3/B sky130_fd_sc_hd__a21o_1_0/a_384_47# 2.82e-20
C221 sky130_fd_sc_hd__xor2_1_3/B sky130_fd_sc_hd__a21o_1_1/a_384_47# 1.76e-19
C222 CI sky130_fd_sc_hd__a21o_1_0/a_81_21# 0.0177f
C223 VPB sky130_fd_sc_hd__xor2_1_3/B 0.167f
C224 S3 sky130_fd_sc_hd__xor2_1_1/a_117_297# 1.88e-20
C225 sky130_fd_sc_hd__xor2_1_1/a_285_297# S1 0.00137f
C226 SUB G2 0.0237f
C227 sky130_fd_sc_hd__a21o_1_0/a_384_47# sky130_fd_sc_hd__xor2_1_2/B 1.35e-20
C228 P1 sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.0139f
C229 P2 G2 6.94e-19
C230 sky130_fd_sc_hd__a21o_1_1/a_384_47# sky130_fd_sc_hd__xor2_1_2/B 4.32e-19
C231 VPB sky130_fd_sc_hd__xor2_1_2/B 0.108f
C232 S2 SUB -0.00162f
C233 P2 S2 0.0068f
C234 sky130_fd_sc_hd__xor2_1_2/a_35_297# S1 2.99e-20
C235 VPB S3 0.041f
C236 sky130_fd_sc_hd__a21o_1_0/a_299_297# VPB 0.0016f
C237 P1 sky130_fd_sc_hd__a21o_1_0/a_384_47# 5.49e-19
C238 sky130_fd_sc_hd__xor2_1_3/B G2 2.64e-19
C239 CI sky130_fd_sc_hd__a21o_1_1/a_81_21# 1.09e-19
C240 sky130_fd_sc_hd__xor2_1_2/a_285_297# S1 4.46e-20
C241 S4 P3 8.8e-19
C242 CI G1 0.0805f
C243 VPB P1 0.00988f
C244 sky130_fd_sc_hd__xor2_1_3/B S2 0.0546f
C245 G1 sky130_fd_sc_hd__a21o_1_0/a_81_21# 0.0272f
C246 G2 sky130_fd_sc_hd__xor2_1_2/B 0.0266f
C247 sky130_fd_sc_hd__xor2_1_2/a_117_297# SUB -0.00177f
C248 sky130_fd_sc_hd__xor2_1_0/a_285_47# SUB -4.65e-19
C249 sky130_fd_sc_hd__xor2_1_0/a_285_47# P2 4.62e-19
C250 sky130_fd_sc_hd__xor2_1_3/a_35_297# SUB 0.00517f
C251 sky130_fd_sc_hd__xor2_1_3/a_35_297# P2 3.67e-21
C252 sky130_fd_sc_hd__xor2_1_1/B S1 0.112f
C253 sky130_fd_sc_hd__xor2_1_1/a_35_297# SUB -0.0109f
C254 S2 sky130_fd_sc_hd__xor2_1_2/B 0.00962f
C255 P2 sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.0178f
C256 sky130_fd_sc_hd__xor2_1_1/B P4 9.9e-21
C257 sky130_fd_sc_hd__xor2_1_0/a_117_297# S1 4.28e-19
C258 VPB sky130_fd_sc_hd__xor2_1_1/a_285_297# 2.35e-20
C259 P1 G2 0.0104f
C260 sky130_fd_sc_hd__a21o_1_2/a_384_47# SUB -2.27e-19
C261 sky130_fd_sc_hd__xor2_1_2/a_117_297# sky130_fd_sc_hd__xor2_1_3/B 0.00134f
C262 S3 S2 0.0102f
C263 sky130_fd_sc_hd__xor2_1_0/a_285_47# sky130_fd_sc_hd__xor2_1_3/B 0.00255f
C264 sky130_fd_sc_hd__xor2_1_3/a_35_297# sky130_fd_sc_hd__xor2_1_3/B 0.0593f
C265 sky130_fd_sc_hd__xor2_1_3/B sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.0714f
C266 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__xor2_1_0/a_285_297# 0.036f
C267 sky130_fd_sc_hd__xor2_1_2/a_117_297# sky130_fd_sc_hd__xor2_1_2/B 0.00267f
C268 VPB sky130_fd_sc_hd__xor2_1_2/a_35_297# 0.00796f
C269 sky130_fd_sc_hd__a21o_1_2/a_384_47# sky130_fd_sc_hd__xor2_1_3/B 0.00131f
C270 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.0678f
C271 sky130_fd_sc_hd__xor2_1_1/B sky130_fd_sc_hd__xor2_1_1/a_117_297# 0.00269f
C272 G3 SUB 8.34e-19
C273 S3 0 0.0366f
C274 P3 0 0.733f
C275 sky130_fd_sc_hd__xor2_1_2/a_285_297# 0 0.00137f
C276 sky130_fd_sc_hd__xor2_1_2/a_35_297# 0 0.255f
C277 SUB 0 1.99f
C278 S2 0 0.0353f
C279 P2 0 0.625f
C280 sky130_fd_sc_hd__xor2_1_1/B 0 0.486f
C281 VPB 0 6.64f
C282 sky130_fd_sc_hd__xor2_1_1/a_285_297# 0 0.00137f
C283 sky130_fd_sc_hd__xor2_1_1/a_35_297# 0 0.255f
C284 S1 0 0.0372f
C285 P1 0 0.561f
C286 CI 0 0.811f
C287 sky130_fd_sc_hd__xor2_1_0/a_285_297# 0 0.00137f
C288 sky130_fd_sc_hd__xor2_1_0/a_35_297# 0 0.255f
C289 sky130_fd_sc_hd__xor2_1_3/B 0 0.336f
C290 sky130_fd_sc_hd__xor2_1_2/B 0 1.53f
C291 G3 0 0.135f
C292 sky130_fd_sc_hd__a21o_1_2/a_299_297# 0 0.0348f
C293 sky130_fd_sc_hd__a21o_1_2/a_81_21# 0 0.147f
C294 G2 0 0.134f
C295 sky130_fd_sc_hd__a21o_1_1/a_299_297# 0 0.0348f
C296 sky130_fd_sc_hd__a21o_1_1/a_81_21# 0 0.147f
C297 G1 0 0.156f
C298 sky130_fd_sc_hd__a21o_1_0/a_299_297# 0 0.0348f
C299 sky130_fd_sc_hd__a21o_1_0/a_81_21# 0 0.147f
C300 S4 0 0.113f
C301 P4 0 0.21f
C302 sky130_fd_sc_hd__xor2_1_3/a_285_297# 0 0.00137f
C303 sky130_fd_sc_hd__xor2_1_3/a_35_297# 0 0.255f
.ends

.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X a_145_75# a_59_75#
X0 VPWR B a_59_75# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.103 pd=0.954 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=6662,278
X1 X a_59_75# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.245 ps=2.27 w=1 l=0.15
**devattr s=6662,278 d=19000,590
X2 VGND B a_145_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0878 pd=0.816 as=0.0567 ps=0.69 w=0.42 l=0.15
**devattr s=2268,138 d=4472,208
X3 a_59_75# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.103 ps=0.954 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
X4 X a_59_75# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.136 ps=1.26 w=0.65 l=0.15
**devattr s=4472,208 d=7280,372
X5 a_145_75# A a_59_75# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.118 ps=1.4 w=0.42 l=0.15
**devattr s=4704,280 d=2268,138
C0 a_59_75# VPWR 0.15f
C1 X B 0.00276f
C2 X VPB 0.0127f
C3 a_145_75# X 5.76e-19
C4 A B 0.0971f
C5 A VPB 0.0806f
C6 VGND B 0.0115f
C7 VGND VPB 0.008f
C8 a_145_75# VGND 0.00468f
C9 A X 1.68e-19
C10 VGND X 0.0993f
C11 VPWR B 0.0117f
C12 VPWR VPB 0.0729f
C13 a_145_75# VPWR 6.31e-19
C14 a_59_75# B 0.143f
C15 a_59_75# VPB 0.0563f
C16 a_59_75# a_145_75# 0.00658f
C17 VPWR X 0.111f
C18 a_59_75# X 0.109f
C19 A VGND 0.0147f
C20 A VPWR 0.0362f
C21 VGND VPWR 0.0461f
C22 A a_59_75# 0.0809f
C23 a_59_75# VGND 0.116f
C24 B VPB 0.0629f
C25 VGND VNB 0.311f
C26 X VNB 0.1f
C27 B VNB 0.113f
C28 A VNB 0.174f
C29 VPWR VNB 0.273f
C30 VPB VNB 0.516f
C31 a_59_75# VNB 0.177f
.ends

.subckt adder_1 A1 B1 A2 B2 A3 B3 A4 B4 G1 P1 G2 P2 G3 P3 G4 P4 sky130_fd_sc_hd__xor2_1_3/a_117_297#
+ sky130_fd_sc_hd__xor2_1_3/a_35_297# sky130_fd_sc_hd__xor2_1_3/a_285_47# sky130_fd_sc_hd__and2_1_3/a_145_75#
+ sky130_fd_sc_hd__and2_1_2/a_59_75# sky130_fd_sc_hd__xor2_1_0/a_285_297# sky130_fd_sc_hd__xor2_1_1/a_285_297#
+ sky130_fd_sc_hd__xor2_1_0/a_35_297# sky130_fd_sc_hd__xor2_1_0/a_285_47# sky130_fd_sc_hd__xor2_1_2/a_285_297#
+ sky130_fd_sc_hd__and2_1_0/a_145_75# sky130_fd_sc_hd__xor2_1_3/a_285_297# sky130_fd_sc_hd__and2_1_3/a_59_75#
+ sky130_fd_sc_hd__xor2_1_1/a_35_297# sky130_fd_sc_hd__xor2_1_1/a_285_47# sky130_fd_sc_hd__and2_1_0/a_59_75#
+ sky130_fd_sc_hd__and2_1_1/a_145_75# sky130_fd_sc_hd__xor2_1_0/a_117_297# sky130_fd_sc_hd__xor2_1_2/a_35_297#
+ sky130_fd_sc_hd__xor2_1_1/a_117_297# sky130_fd_sc_hd__xor2_1_2/a_285_47# sky130_fd_sc_hd__and2_1_2/a_145_75#
+ SUB sky130_fd_sc_hd__and2_1_1/a_59_75# sky130_fd_sc_hd__xor2_1_2/a_117_297# VDD
Xsky130_fd_sc_hd__xor2_1_3 A4 B4 SUB SUB VDD VDD P4 sky130_fd_sc_hd__xor2_1_3/a_117_297#
+ sky130_fd_sc_hd__xor2_1_3/a_285_297# sky130_fd_sc_hd__xor2_1_3/a_285_47# sky130_fd_sc_hd__xor2_1_3/a_35_297#
+ sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__and2_1_0 A1 B1 SUB SUB VDD VDD G1 sky130_fd_sc_hd__and2_1_0/a_145_75#
+ sky130_fd_sc_hd__and2_1_0/a_59_75# sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__and2_1_1 A2 B2 SUB SUB VDD VDD G2 sky130_fd_sc_hd__and2_1_1/a_145_75#
+ sky130_fd_sc_hd__and2_1_1/a_59_75# sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__and2_1_2 A3 B3 SUB SUB VDD VDD G3 sky130_fd_sc_hd__and2_1_2/a_145_75#
+ sky130_fd_sc_hd__and2_1_2/a_59_75# sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__and2_1_3 A4 B4 SUB SUB VDD VDD G4 sky130_fd_sc_hd__and2_1_3/a_145_75#
+ sky130_fd_sc_hd__and2_1_3/a_59_75# sky130_fd_sc_hd__and2_1
Xsky130_fd_sc_hd__xor2_1_0 A1 B1 SUB SUB VDD VDD P1 sky130_fd_sc_hd__xor2_1_0/a_117_297#
+ sky130_fd_sc_hd__xor2_1_0/a_285_297# sky130_fd_sc_hd__xor2_1_0/a_285_47# sky130_fd_sc_hd__xor2_1_0/a_35_297#
+ sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_1 A2 B2 SUB SUB VDD VDD P2 sky130_fd_sc_hd__xor2_1_1/a_117_297#
+ sky130_fd_sc_hd__xor2_1_1/a_285_297# sky130_fd_sc_hd__xor2_1_1/a_285_47# sky130_fd_sc_hd__xor2_1_1/a_35_297#
+ sky130_fd_sc_hd__xor2_1
Xsky130_fd_sc_hd__xor2_1_2 A3 B3 SUB SUB VDD VDD P3 sky130_fd_sc_hd__xor2_1_2/a_117_297#
+ sky130_fd_sc_hd__xor2_1_2/a_285_297# sky130_fd_sc_hd__xor2_1_2/a_285_47# sky130_fd_sc_hd__xor2_1_2/a_35_297#
+ sky130_fd_sc_hd__xor2_1
C0 P3 sky130_fd_sc_hd__xor2_1_3/a_285_297# 9.07e-20
C1 G2 G3 -1.94e-25
C2 A1 B2 1.47e-19
C3 A4 B4 0.249f
C4 B4 sky130_fd_sc_hd__xor2_1_3/a_285_47# 2.19e-19
C5 A4 G3 1.39e-19
C6 G4 sky130_fd_sc_hd__xor2_1_3/a_285_297# 6.56e-19
C7 P1 A2 0.0305f
C8 sky130_fd_sc_hd__and2_1_3/a_59_75# sky130_fd_sc_hd__xor2_1_2/a_35_297# 0.00179f
C9 sky130_fd_sc_hd__and2_1_2/a_59_75# sky130_fd_sc_hd__xor2_1_2/a_35_297# 5.6e-19
C10 sky130_fd_sc_hd__xor2_1_2/a_35_297# B3 0.0715f
C11 sky130_fd_sc_hd__xor2_1_2/a_35_297# P4 5.81e-21
C12 SUB P1 0.0117f
C13 G1 sky130_fd_sc_hd__xor2_1_0/a_285_297# 5.75e-19
C14 A2 sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.0397f
C15 sky130_fd_sc_hd__xor2_1_0/a_117_297# SUB -0.00177f
C16 sky130_fd_sc_hd__xor2_1_2/a_285_297# VDD 4.65e-20
C17 B4 sky130_fd_sc_hd__xor2_1_2/a_35_297# 4.2e-19
C18 G3 sky130_fd_sc_hd__xor2_1_2/a_35_297# 0.0665f
C19 B1 sky130_fd_sc_hd__xor2_1_0/a_285_297# 1.19e-19
C20 SUB sky130_fd_sc_hd__xor2_1_1/a_35_297# -0.00565f
C21 sky130_fd_sc_hd__and2_1_3/a_59_75# P3 0.00722f
C22 sky130_fd_sc_hd__and2_1_2/a_59_75# P3 9.47e-20
C23 B3 P3 0.00724f
C24 P4 P3 2.91e-20
C25 P1 P2 3.79e-19
C26 sky130_fd_sc_hd__and2_1_3/a_59_75# G4 0.0026f
C27 sky130_fd_sc_hd__xor2_1_0/a_35_297# G1 0.0663f
C28 G4 B3 9.35e-20
C29 B4 P3 7.42e-19
C30 G4 P4 0.00346f
C31 P1 sky130_fd_sc_hd__and2_1_1/a_59_75# 0.00746f
C32 B1 G1 0.0397f
C33 G3 P3 2.77e-19
C34 B1 sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.0359f
C35 sky130_fd_sc_hd__xor2_1_1/a_35_297# P2 0.00234f
C36 G4 B4 0.0423f
C37 B3 sky130_fd_sc_hd__and2_1_2/a_145_75# 2.46e-20
C38 sky130_fd_sc_hd__and2_1_1/a_59_75# sky130_fd_sc_hd__xor2_1_1/a_35_297# 5.6e-19
C39 G2 P1 6.62e-19
C40 P4 sky130_fd_sc_hd__xor2_1_3/a_285_297# 0.0109f
C41 sky130_fd_sc_hd__xor2_1_0/a_117_297# G2 1.14e-19
C42 G4 G3 0.00197f
C43 sky130_fd_sc_hd__xor2_1_1/a_285_47# B2 2.25e-19
C44 A2 VDD 0.198f
C45 B4 sky130_fd_sc_hd__xor2_1_3/a_285_297# 1.19e-19
C46 G2 sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.0663f
C47 sky130_fd_sc_hd__xor2_1_1/a_285_297# A2 6.41e-19
C48 P1 sky130_fd_sc_hd__xor2_1_1/a_117_297# 1.21e-19
C49 SUB VDD -0.222f
C50 sky130_fd_sc_hd__and2_1_0/a_145_75# VDD -6.31e-19
C51 B2 A2 0.256f
C52 sky130_fd_sc_hd__and2_1_3/a_59_75# B3 4.1e-19
C53 sky130_fd_sc_hd__and2_1_2/a_59_75# B3 0.0565f
C54 A3 sky130_fd_sc_hd__xor2_1_2/a_285_297# 6.24e-19
C55 sky130_fd_sc_hd__and2_1_3/a_59_75# P4 2.68e-20
C56 SUB B2 0.157f
C57 sky130_fd_sc_hd__and2_1_0/a_59_75# G1 0.00228f
C58 sky130_fd_sc_hd__xor2_1_2/a_117_297# VDD -1.39e-19
C59 sky130_fd_sc_hd__and2_1_0/a_59_75# sky130_fd_sc_hd__xor2_1_0/a_35_297# 5.6e-19
C60 P2 VDD 0.0747f
C61 sky130_fd_sc_hd__and2_1_0/a_145_75# B2 1.12e-21
C62 sky130_fd_sc_hd__and2_1_3/a_59_75# B4 0.0576f
C63 B4 B3 0.00433f
C64 sky130_fd_sc_hd__xor2_1_3/a_117_297# VDD -1.39e-19
C65 sky130_fd_sc_hd__xor2_1_1/a_285_297# P2 0.0109f
C66 sky130_fd_sc_hd__and2_1_1/a_59_75# VDD -7.45e-19
C67 sky130_fd_sc_hd__and2_1_0/a_59_75# B1 0.0544f
C68 sky130_fd_sc_hd__and2_1_3/a_59_75# G3 9.08e-20
C69 B4 P4 0.00126f
C70 sky130_fd_sc_hd__and2_1_2/a_59_75# G3 0.0029f
C71 G3 B3 0.0409f
C72 G2 VDD 0.0388f
C73 B2 P2 0.00129f
C74 G2 sky130_fd_sc_hd__xor2_1_1/a_285_297# 5.75e-19
C75 B4 G3 3.51e-20
C76 P3 sky130_fd_sc_hd__xor2_1_1/a_35_297# 1.16e-20
C77 A4 VDD 0.197f
C78 sky130_fd_sc_hd__and2_1_1/a_59_75# B2 0.0564f
C79 P1 sky130_fd_sc_hd__xor2_1_0/a_285_297# 0.00448f
C80 SUB sky130_fd_sc_hd__xor2_1_2/a_285_47# -2.55e-19
C81 G2 B2 0.042f
C82 A3 A2 0.00809f
C83 sky130_fd_sc_hd__xor2_1_1/a_117_297# VDD -1.39e-19
C84 P1 G1 3.4e-19
C85 A3 SUB 0.0164f
C86 sky130_fd_sc_hd__xor2_1_0/a_117_297# G1 7.26e-19
C87 P1 sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.00153f
C88 sky130_fd_sc_hd__xor2_1_2/a_35_297# VDD 0.0079f
C89 sky130_fd_sc_hd__xor2_1_0/a_285_47# B2 5.6e-20
C90 B1 P1 0.0021f
C91 A1 A2 0.00698f
C92 SUB sky130_fd_sc_hd__xor2_1_3/a_35_297# -0.0066f
C93 sky130_fd_sc_hd__xor2_1_2/a_117_297# A3 0.00414f
C94 A3 P2 0.00732f
C95 SUB A1 0.0438f
C96 P3 VDD 0.0448f
C97 A3 sky130_fd_sc_hd__and2_1_1/a_59_75# 3.22e-20
C98 sky130_fd_sc_hd__and2_1_0/a_145_75# A1 0.00119f
C99 sky130_fd_sc_hd__xor2_1_1/a_285_297# P3 2.3e-20
C100 sky130_fd_sc_hd__and2_1_2/a_59_75# sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.00133f
C101 B3 sky130_fd_sc_hd__xor2_1_1/a_35_297# 4e-19
C102 G4 VDD 0.0395f
C103 G2 A3 6.19e-20
C104 sky130_fd_sc_hd__xor2_1_0/a_285_297# VDD 4.65e-20
C105 A4 A3 0.00249f
C106 A1 P2 1.59e-21
C107 sky130_fd_sc_hd__xor2_1_3/a_285_297# VDD 3.2e-32
C108 sky130_fd_sc_hd__and2_1_2/a_145_75# VDD -6.31e-19
C109 sky130_fd_sc_hd__and2_1_0/a_59_75# P1 1.33e-19
C110 G1 VDD 0.0385f
C111 sky130_fd_sc_hd__xor2_1_0/a_35_297# VDD 0.00867f
C112 A4 sky130_fd_sc_hd__xor2_1_3/a_35_297# 0.0402f
C113 G2 A1 1.14e-19
C114 B1 VDD 0.00679f
C115 B2 sky130_fd_sc_hd__and2_1_2/a_145_75# 2.37e-21
C116 SUB sky130_fd_sc_hd__xor2_1_2/a_285_297# -0.00166f
C117 A3 sky130_fd_sc_hd__xor2_1_2/a_35_297# 0.0336f
C118 G1 B2 7.99e-20
C119 sky130_fd_sc_hd__xor2_1_0/a_35_297# B2 7.19e-19
C120 A4 sky130_fd_sc_hd__and2_1_3/a_145_75# 0.00119f
C121 sky130_fd_sc_hd__and2_1_3/a_59_75# VDD -7.45e-19
C122 sky130_fd_sc_hd__and2_1_2/a_59_75# VDD 0.00479f
C123 B3 VDD 0.0264f
C124 B1 B2 0.00218f
C125 P4 VDD 0.0238f
C126 sky130_fd_sc_hd__xor2_1_2/a_285_297# P2 2.5e-20
C127 A3 P3 0.006f
C128 B4 VDD 0.00646f
C129 sky130_fd_sc_hd__and2_1_2/a_59_75# B2 1.27e-19
C130 B3 B2 0.00271f
C131 G3 VDD 0.0413f
C132 A3 G4 1.26e-19
C133 sky130_fd_sc_hd__xor2_1_0/a_117_297# P1 3.4e-19
C134 P3 sky130_fd_sc_hd__xor2_1_3/a_35_297# 1.05e-19
C135 SUB A2 0.0431f
C136 A4 sky130_fd_sc_hd__xor2_1_2/a_285_297# 3.31e-19
C137 P1 sky130_fd_sc_hd__xor2_1_1/a_35_297# 1.51e-19
C138 sky130_fd_sc_hd__and2_1_0/a_59_75# VDD -0.00241f
C139 A3 sky130_fd_sc_hd__and2_1_2/a_145_75# 0.00119f
C140 G4 sky130_fd_sc_hd__xor2_1_3/a_35_297# 0.0665f
C141 A1 sky130_fd_sc_hd__xor2_1_0/a_285_297# 6.41e-19
C142 sky130_fd_sc_hd__and2_1_1/a_145_75# VDD -6.31e-19
C143 sky130_fd_sc_hd__and2_1_0/a_59_75# B2 5.54e-20
C144 A2 P2 0.00233f
C145 B3 sky130_fd_sc_hd__xor2_1_2/a_285_47# 0.00257f
C146 sky130_fd_sc_hd__and2_1_1/a_59_75# A2 0.0589f
C147 sky130_fd_sc_hd__xor2_1_2/a_117_297# SUB -0.00177f
C148 SUB P2 0.00985f
C149 sky130_fd_sc_hd__and2_1_1/a_145_75# B2 2.28e-20
C150 A3 sky130_fd_sc_hd__and2_1_2/a_59_75# 0.0594f
C151 G1 A1 0.0701f
C152 SUB sky130_fd_sc_hd__xor2_1_3/a_117_297# -0.00177f
C153 A3 B3 0.294f
C154 G2 A2 0.071f
C155 SUB sky130_fd_sc_hd__and2_1_1/a_59_75# 0.00649f
C156 sky130_fd_sc_hd__xor2_1_0/a_35_297# A1 0.0402f
C157 A3 P4 3.19e-21
C158 B1 A1 0.264f
C159 G2 SUB -1.95e-19
C160 sky130_fd_sc_hd__xor2_1_2/a_285_297# P3 0.00179f
C161 P1 VDD 0.0465f
C162 sky130_fd_sc_hd__xor2_1_2/a_117_297# P2 1.97e-20
C163 sky130_fd_sc_hd__xor2_1_0/a_117_297# VDD -1.39e-19
C164 sky130_fd_sc_hd__and2_1_3/a_59_75# sky130_fd_sc_hd__xor2_1_3/a_35_297# 5.6e-19
C165 A3 G3 0.074f
C166 A4 SUB 0.0446f
C167 P1 sky130_fd_sc_hd__xor2_1_1/a_285_297# 1.46e-19
C168 sky130_fd_sc_hd__xor2_1_1/a_117_297# A2 0.00414f
C169 P4 sky130_fd_sc_hd__xor2_1_3/a_35_297# 0.00234f
C170 sky130_fd_sc_hd__and2_1_1/a_59_75# P2 4.05e-20
C171 G4 sky130_fd_sc_hd__xor2_1_2/a_285_297# 3.71e-19
C172 sky130_fd_sc_hd__xor2_1_1/a_35_297# VDD 0.00949f
C173 P1 B2 8.23e-19
C174 SUB sky130_fd_sc_hd__xor2_1_1/a_117_297# -0.00177f
C175 B4 sky130_fd_sc_hd__xor2_1_3/a_35_297# 0.0414f
C176 G2 P2 0.00318f
C177 G3 sky130_fd_sc_hd__xor2_1_3/a_35_297# 5.99e-22
C178 B3 sky130_fd_sc_hd__and2_1_3/a_145_75# 6.15e-21
C179 G2 sky130_fd_sc_hd__and2_1_1/a_59_75# 0.00228f
C180 B2 sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.0446f
C181 A4 sky130_fd_sc_hd__xor2_1_3/a_117_297# 0.00414f
C182 SUB sky130_fd_sc_hd__xor2_1_2/a_35_297# -0.0109f
C183 sky130_fd_sc_hd__xor2_1_1/a_117_297# P2 5.63e-19
C184 B4 sky130_fd_sc_hd__and2_1_3/a_145_75# 2.46e-20
C185 sky130_fd_sc_hd__and2_1_0/a_59_75# A1 0.0581f
C186 SUB P3 0.0125f
C187 sky130_fd_sc_hd__xor2_1_2/a_35_297# P2 1.96e-20
C188 G2 sky130_fd_sc_hd__xor2_1_1/a_117_297# 7.26e-19
C189 sky130_fd_sc_hd__xor2_1_0/a_285_297# A2 3.31e-19
C190 sky130_fd_sc_hd__xor2_1_2/a_285_297# B3 0.00523f
C191 sky130_fd_sc_hd__xor2_1_2/a_285_297# P4 2.02e-20
C192 G4 SUB -1.95e-19
C193 sky130_fd_sc_hd__xor2_1_1/a_285_297# VDD 6.02e-20
C194 A3 P1 1.12e-21
C195 sky130_fd_sc_hd__xor2_1_2/a_117_297# P3 2.16e-19
C196 P3 P2 2.24e-20
C197 G1 A2 1.33e-19
C198 sky130_fd_sc_hd__xor2_1_2/a_285_297# G3 6.58e-19
C199 B2 VDD 0.00698f
C200 A4 sky130_fd_sc_hd__xor2_1_2/a_35_297# 0.0101f
C201 sky130_fd_sc_hd__xor2_1_0/a_35_297# A2 0.0101f
C202 A3 sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.00595f
C203 sky130_fd_sc_hd__xor2_1_3/a_117_297# P3 7.54e-20
C204 sky130_fd_sc_hd__xor2_1_1/a_285_47# B3 3.82e-20
C205 sky130_fd_sc_hd__xor2_1_1/a_285_297# B2 1.19e-19
C206 sky130_fd_sc_hd__xor2_1_2/a_117_297# G4 1.25e-19
C207 B1 A2 0.00281f
C208 SUB G1 0.00116f
C209 SUB sky130_fd_sc_hd__xor2_1_0/a_35_297# -0.00339f
C210 sky130_fd_sc_hd__xor2_1_0/a_285_297# P2 1.01e-20
C211 G4 sky130_fd_sc_hd__xor2_1_3/a_117_297# 7.98e-19
C212 P1 A1 0.00719f
C213 sky130_fd_sc_hd__xor2_1_0/a_117_297# A1 0.00414f
C214 B1 SUB 0.134f
C215 A4 P3 0.0296f
C216 B3 A2 1e-19
C217 G2 sky130_fd_sc_hd__xor2_1_0/a_285_297# 3.25e-19
C218 A4 G4 0.0729f
C219 sky130_fd_sc_hd__xor2_1_0/a_35_297# P2 2.9e-21
C220 sky130_fd_sc_hd__and2_1_3/a_59_75# SUB 0.00649f
C221 SUB sky130_fd_sc_hd__and2_1_2/a_59_75# 0.00617f
C222 sky130_fd_sc_hd__xor2_1_2/a_285_47# VDD -8.2e-19
C223 SUB B3 0.232f
C224 sky130_fd_sc_hd__and2_1_1/a_59_75# G1 8.11e-20
C225 SUB P4 0.00985f
C226 sky130_fd_sc_hd__and2_1_1/a_59_75# sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.00179f
C227 A4 sky130_fd_sc_hd__xor2_1_3/a_285_297# 6.41e-19
C228 B1 sky130_fd_sc_hd__and2_1_1/a_59_75# 9.42e-20
C229 G2 G1 0.00179f
C230 sky130_fd_sc_hd__xor2_1_2/a_35_297# P3 0.00192f
C231 SUB B4 0.154f
C232 A3 VDD 0.208f
C233 G2 sky130_fd_sc_hd__xor2_1_0/a_35_297# 2.05e-19
C234 SUB G3 -1.95e-19
C235 A3 sky130_fd_sc_hd__xor2_1_1/a_285_297# 4.35e-19
C236 sky130_fd_sc_hd__and2_1_2/a_59_75# P2 0.00164f
C237 B3 P2 5.55e-19
C238 sky130_fd_sc_hd__and2_1_0/a_59_75# A2 4.2e-20
C239 G2 B1 8.95e-20
C240 G4 sky130_fd_sc_hd__xor2_1_2/a_35_297# 2.26e-19
C241 P4 sky130_fd_sc_hd__xor2_1_3/a_117_297# 5.63e-19
C242 sky130_fd_sc_hd__and2_1_0/a_59_75# SUB -0.00661f
C243 A3 B2 0.00246f
C244 sky130_fd_sc_hd__xor2_1_3/a_35_297# VDD 0.00289f
C245 sky130_fd_sc_hd__xor2_1_2/a_117_297# G3 7.99e-19
C246 sky130_fd_sc_hd__and2_1_1/a_145_75# A2 0.00119f
C247 G3 P2 0.00384f
C248 A1 VDD 0.182f
C249 B1 sky130_fd_sc_hd__xor2_1_0/a_285_47# 2.19e-19
C250 sky130_fd_sc_hd__and2_1_3/a_59_75# A4 0.0591f
C251 A4 sky130_fd_sc_hd__and2_1_2/a_59_75# 4.2e-20
C252 G3 sky130_fd_sc_hd__xor2_1_3/a_117_297# 9e-22
C253 A4 B3 0.00861f
C254 G4 P3 5.33e-19
C255 A4 P4 0.00232f
C256 sky130_fd_sc_hd__and2_1_3/a_145_75# VDD -6.31e-19
C257 G1 0 0.0305f
C258 SUB 0 2.81f
C259 VDD 0 7.09f
C260 P3 0 0.0173f
C261 sky130_fd_sc_hd__xor2_1_2/a_285_297# 0 0.00137f
C262 sky130_fd_sc_hd__xor2_1_2/a_35_297# 0 0.255f
C263 P2 0 0.0182f
C264 A2 0 0.317f
C265 B2 0 0.338f
C266 sky130_fd_sc_hd__xor2_1_1/a_285_297# 0 0.00137f
C267 sky130_fd_sc_hd__xor2_1_1/a_35_297# 0 0.255f
C268 P1 0 0.0183f
C269 A1 0 0.373f
C270 B1 0 0.337f
C271 sky130_fd_sc_hd__xor2_1_0/a_285_297# 0 0.00137f
C272 sky130_fd_sc_hd__xor2_1_0/a_35_297# 0 0.255f
C273 G4 0 0.0255f
C274 B4 0 0.342f
C275 A4 0 0.328f
C276 sky130_fd_sc_hd__and2_1_3/a_59_75# 0 0.177f
C277 G3 0 0.0256f
C278 B3 0 0.339f
C279 A3 0 0.323f
C280 sky130_fd_sc_hd__and2_1_2/a_59_75# 0 0.177f
C281 G2 0 0.0255f
C282 sky130_fd_sc_hd__and2_1_1/a_59_75# 0 0.177f
C283 sky130_fd_sc_hd__and2_1_0/a_59_75# 0 0.177f
C284 P4 0 0.0763f
C285 sky130_fd_sc_hd__xor2_1_3/a_285_297# 0 0.00137f
C286 sky130_fd_sc_hd__xor2_1_3/a_35_297# 0 0.255f
.ends

.subckt adder_4 A1 B1 A2 B2 A3 B3 A4 B4 CI S1 S2 S3 S4 CO VDD GND
Xadder_2_0 CI adder_3_0/P1 adder_3_0/G1 adder_3_0/P2 adder_3_0/G2 adder_3_0/P3 adder_3_0/G3
+ adder_3_0/P4 adder_2_0/G4 CO adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47#
+ adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_384_47# adder_2_0/sky130_fd_sc_hd__a21o_1_1/X
+ adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_299_297#
+ VDD adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_384_47#
+ adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# adder_2_0/sky130_fd_sc_hd__and4_1_0/a_109_47#
+ adder_2_0/sky130_fd_sc_hd__a21o_1_2/X adder_2_0/sky130_fd_sc_hd__a21o_1_0/X adder_2_0/sky130_fd_sc_hd__and4_1_0/X
+ adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21#
+ GND adder_2_0/sky130_fd_sc_hd__and4_1_0/a_197_47# adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_384_47#
+ adder_2_0/sky130_fd_sc_hd__and4_1_0/a_303_47# adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21#
+ adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_384_47# adder_2
Xadder_3_0 adder_3_0/G1 adder_3_0/P2 adder_3_0/G2 adder_3_0/G3 adder_3_0/P4 S1 S2
+ S3 S4 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_117_297# adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297#
+ adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_47#
+ adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_384_47#
+ adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297#
+ adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_47# adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21#
+ adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297#
+ adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297#
+ adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297#
+ adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_47#
+ adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21#
+ adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297#
+ adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_47# adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_117_297#
+ CI adder_3_0/P1 GND adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_117_297#
+ VDD adder_3_0/P3 adder_3
Xadder_1_0 A1 B1 A2 B2 A3 B3 A4 B4 adder_3_0/G1 adder_3_0/P1 adder_3_0/G2 adder_3_0/P2
+ adder_3_0/G3 adder_3_0/P3 adder_2_0/G4 adder_3_0/P4 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_117_297#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_47#
+ adder_1_0/sky130_fd_sc_hd__and2_1_3/a_145_75# adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_47#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# adder_1_0/sky130_fd_sc_hd__and2_1_0/a_145_75#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_47#
+ adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# adder_1_0/sky130_fd_sc_hd__and2_1_1/a_145_75#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_117_297# adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_47#
+ adder_1_0/sky130_fd_sc_hd__and2_1_2/a_145_75# GND adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75#
+ adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# VDD adder_1
C0 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 0.00297f
C1 adder_3_0/P2 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_47# -4.62e-19
C2 adder_3_0/P2 S3 3.05e-21
C3 B2 GND 0.00396f
C4 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B GND 0.00204f
C5 S4 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_47# 0.00104f
C6 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_3_0/P2 0.00628f
C7 adder_3_0/P2 adder_2_0/G4 0.0231f
C8 A3 VDD 0.208f
C9 S1 adder_2_0/sky130_fd_sc_hd__and4_1_0/X 0.00171f
C10 A3 B3 1.3f
C11 adder_3_0/P3 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 1.67e-19
C12 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_47# VDD -8.51e-21
C13 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_47# B3 5.14e-19
C14 adder_3_0/G3 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_117_297# 8.67e-21
C15 B4 CI 1.51f
C16 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# CI 2.49e-19
C17 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# B2 6.12e-20
C18 adder_3_0/P2 S2 0.0771f
C19 adder_3_0/G3 adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 2.97e-20
C20 adder_3_0/P3 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.00106f
C21 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_3_0/P3 0.011f
C22 adder_3_0/P1 adder_3_0/G2 0.405f
C23 adder_3_0/G3 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 2.64e-19
C24 adder_3_0/P4 adder_3_0/G2 4.99e-20
C25 A3 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_117_297# 2.11e-19
C26 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_145_75# adder_3_0/G1 0.00101f
C27 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 3.16e-19
C28 B1 CI 1.95e-19
C29 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 2.93e-19
C30 CO adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 0.0284f
C31 adder_3_0/P4 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 3.55e-20
C32 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# CI 0.00104f
C33 adder_3_0/P2 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 0.0124f
C34 adder_3_0/P3 adder_1_0/sky130_fd_sc_hd__and2_1_3/a_145_75# 6.88e-19
C35 adder_3_0/P3 A4 0.0462f
C36 adder_2_0/G4 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.00465f
C37 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 7.55e-22
C38 adder_3_0/P4 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_117_297# 9.54e-19
C39 A2 GND 0.00582f
C40 adder_3_0/P3 VDD 0.534f
C41 adder_3_0/G1 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 1.03e-19
C42 adder_3_0/P3 B3 0.0502f
C43 CO adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.00229f
C44 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X GND 1.34e-19
C45 adder_3_0/G3 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# 3.12e-19
C46 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# A4 3.72e-20
C47 adder_2_0/G4 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 7.97e-20
C48 S1 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 3.99e-19
C49 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# A2 0.00125f
C50 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_2_0/G4 1.9e-19
C51 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# VDD 0.00935f
C52 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# B3 4.65e-20
C53 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# GND 7.61e-19
C54 CO adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 0.00806f
C55 adder_3_0/G2 CI 0.0259f
C56 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_3_0/P1 0.00384f
C57 adder_3_0/P2 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.00226f
C58 adder_3_0/P2 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_145_75# 4.99e-19
C59 adder_3_0/P1 B2 0.00166f
C60 adder_3_0/G3 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0.00128f
C61 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_3_0/P1 0.0196f
C62 A1 A4 2.8e-19
C63 adder_3_0/P4 B2 6.88e-19
C64 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_3_0/P4 1.5e-19
C65 CO adder_2_0/sky130_fd_sc_hd__and4_1_0/X 0.106f
C66 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 2.13e-20
C67 adder_2_0/G4 adder_1_0/sky130_fd_sc_hd__and2_1_3/a_145_75# 8.23e-19
C68 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# GND 1.54e-19
C69 VDD A1 0.37f
C70 adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# adder_3_0/P3 0.00388f
C71 adder_2_0/G4 A4 0.0821f
C72 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# CI 5.48e-19
C73 A1 B3 3.87e-19
C74 VDD S3 8.27e-19
C75 adder_3_0/P2 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 0.0148f
C76 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B VDD -2.88e-19
C77 adder_2_0/G4 VDD 0.174f
C78 adder_2_0/G4 B3 2.86e-19
C79 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_3_0/P2 -9.82e-21
C80 S4 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# -1.86e-19
C81 adder_2_0/sky130_fd_sc_hd__and4_1_0/X GND 1.11e-19
C82 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# adder_3_0/P3 0.00405f
C83 adder_3_0/P4 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_47# 5.65e-19
C84 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# adder_3_0/P3 0.00147f
C85 S4 S1 0.0283f
C86 CO S1 0.257f
C87 VDD S2 0.00253f
C88 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 2.45e-19
C89 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# S1 1.21e-20
C90 adder_3_0/G3 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.0147f
C91 adder_3_0/G3 B4 9.64e-20
C92 CO adder_2_0/sky130_fd_sc_hd__and4_1_0/a_109_47# 3.18e-19
C93 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# GND 8.85e-19
C94 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_3_0/sky130_fd_sc_hd__xor2_1_2/B -9.88e-19
C95 adder_3_0/P2 A4 1.08e-19
C96 adder_3_0/G3 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 0.00432f
C97 S1 GND 1.14f
C98 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# CI 3.01e-20
C99 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 9.14e-21
C100 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# adder_3_0/sky130_fd_sc_hd__xor2_1_2/B -2.17e-19
C101 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# adder_3_0/sky130_fd_sc_hd__xor2_1_2/B -7.49e-19
C102 adder_3_0/P2 VDD 0.267f
C103 B2 CI 3.41e-19
C104 adder_3_0/P2 B3 8.59e-19
C105 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B CI 0.0245f
C106 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_2_0/sky130_fd_sc_hd__and4_1_0/X 1.35e-19
C107 adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# adder_2_0/G4 0.0161f
C108 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X adder_2_0/sky130_fd_sc_hd__a21o_1_1/X -9.62e-21
C109 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_384_47# CO 3.28e-19
C110 GND adder_2_0/sky130_fd_sc_hd__a21o_1_1/X -6.74e-19
C111 A2 adder_3_0/P1 0.0449f
C112 adder_3_0/P4 A2 4.36e-19
C113 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# GND 9.8e-19
C114 B4 A3 8.32e-19
C115 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# VDD 6.51e-19
C116 VDD adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 5.68e-32
C117 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X adder_3_0/P1 0.0274f
C118 adder_3_0/P4 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 0.0226f
C119 adder_3_0/G3 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_145_75# 1.86e-19
C120 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X adder_3_0/G1 0.0445f
C121 B1 adder_3_0/G3 0.00439f
C122 adder_3_0/G1 GND 0.376f
C123 S4 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 0.0084f
C124 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# adder_3_0/G1 0.0118f
C125 CO adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 2.53e-19
C126 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# adder_2_0/G4 1.65e-19
C127 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 5.31e-21
C128 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# adder_2_0/G4 0.00559f
C129 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_3_0/P1 7.47e-19
C130 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# CI 0.00225f
C131 adder_3_0/P4 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_47# 0.00104f
C132 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# S1 -0.00115f
C133 adder_3_0/P4 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 3.44e-19
C134 adder_2_0/sky130_fd_sc_hd__and4_1_0/X adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 5.71e-20
C135 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_3_0/G1 0.00976f
C136 adder_3_0/P2 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_117_297# 0.00103f
C137 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# adder_3_0/P3 0.0039f
C138 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# GND 0.00127f
C139 B1 A3 9.01e-19
C140 adder_3_0/P3 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 4.09e-20
C141 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_2_0/sky130_fd_sc_hd__a21o_1_1/X -4.9e-21
C142 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# adder_3_0/P1 0.0174f
C143 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# S1 -6.35e-20
C144 adder_3_0/P4 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# -2.26e-19
C145 VDD adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.00242f
C146 S1 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# -7.29e-19
C147 adder_3_0/P2 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# -1.11e-20
C148 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 3.33e-20
C149 adder_3_0/G3 adder_3_0/G2 0.882f
C150 A2 CI 2.43e-19
C151 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# A4 6.49e-20
C152 adder_2_0/sky130_fd_sc_hd__and4_1_0/X adder_3_0/P1 0.00468f
C153 adder_3_0/P4 adder_2_0/sky130_fd_sc_hd__and4_1_0/X 2.22e-19
C154 adder_3_0/G2 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.0946f
C155 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X CI 0.0104f
C156 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# A4 0.00128f
C157 adder_3_0/P3 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.00509f
C158 B4 adder_3_0/P3 0.00132f
C159 S4 CO 0.209f
C160 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# VDD -6.01e-19
C161 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# B3 2.25e-20
C162 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# CO 0.00874f
C163 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# VDD -6.68e-19
C164 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# B3 0.0107f
C165 adder_3_0/G3 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 0.0163f
C166 adder_3_0/P3 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# 0.00275f
C167 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# adder_3_0/P3 0.0383f
C168 adder_3_0/G3 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_117_297# -9e-22
C169 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# CI 3.33e-19
C170 adder_3_0/P4 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 0.0141f
C171 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# B4 3.05e-20
C172 S4 GND 0.0982f
C173 A3 adder_3_0/G2 2.08e-19
C174 adder_3_0/G3 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_384_47# 4.39e-19
C175 CO GND 0.151f
C176 S1 adder_3_0/P1 0.0451f
C177 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# GND 1.4e-19
C178 adder_3_0/P4 S1 0.00107f
C179 adder_2_0/G4 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 2.44e-19
C180 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_384_47# adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 7.63e-20
C181 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 2.84e-20
C182 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# GND 4.55e-19
C183 adder_3_0/P1 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 0.0208f
C184 VDD A4 0.142f
C185 adder_3_0/P4 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 0.00539f
C186 A3 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 0.0163f
C187 A4 B3 1.7f
C188 adder_3_0/P4 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 0.0131f
C189 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X GND 6.92e-20
C190 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# CI 0.00244f
C191 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# adder_3_0/G1 0.00311f
C192 VDD B3 0.171f
C193 adder_3_0/P1 adder_3_0/G1 0.0488f
C194 B4 A1 2.13e-19
C195 adder_3_0/P4 adder_3_0/G1 1.36e-20
C196 B1 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# 6.38e-19
C197 adder_3_0/G3 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 0.00261f
C198 B4 adder_2_0/G4 0.0886f
C199 adder_2_0/G4 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.00122f
C200 adder_2_0/sky130_fd_sc_hd__and4_1_0/X CI 0.0231f
C201 adder_3_0/P2 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 1.63e-19
C202 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 8.3e-19
C203 adder_3_0/P2 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# -1.01e-20
C204 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# GND -5.32e-19
C205 adder_3_0/G3 B2 0.00108f
C206 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_3_0/G3 0.0318f
C207 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# CO 0.014f
C208 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 6.98e-20
C209 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# 4.05e-20
C210 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# adder_2_0/G4 9.53e-20
C211 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_3_0/sky130_fd_sc_hd__xor2_1_2/B -0.014f
C212 adder_3_0/P4 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 0.00776f
C213 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 0.00285f
C214 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_384_47# adder_3_0/G1 4.44e-19
C215 adder_3_0/P1 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 1.34e-20
C216 B1 A1 0.237f
C217 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# GND 8.68e-19
C218 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# A3 5.96e-20
C219 adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# A4 0.0161f
C220 S1 CI 4.68e-19
C221 adder_3_0/P3 adder_3_0/G2 0.0027f
C222 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# GND 9.7e-20
C223 A3 B2 0.938f
C224 adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# VDD -5.1e-20
C225 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# A1 9.74e-19
C226 adder_3_0/G3 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# 3.28e-19
C227 CO adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 0.00441f
C228 B4 adder_3_0/P2 9.02e-20
C229 adder_3_0/P2 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.00106f
C230 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_109_47# CI 3.82e-20
C231 CI adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 2.11e-19
C232 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# A4 0.00264f
C233 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# S1 -3.09e-20
C234 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 1.46e-20
C235 adder_3_0/P3 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 7.39e-20
C236 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 2.6e-20
C237 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# adder_3_0/G2 7.89e-19
C238 adder_3_0/P2 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# 2.5e-19
C239 adder_3_0/G1 CI 0.0965f
C240 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# B3 0.0195f
C241 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_117_297# adder_3_0/P3 3.36e-20
C242 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_384_47# CI 6.1e-19
C243 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_384_47# adder_3_0/P3 4.84e-19
C244 adder_3_0/G3 A2 0.0115f
C245 adder_3_0/P4 S4 0.0312f
C246 CO adder_3_0/P1 0.0294f
C247 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# adder_3_0/P1 0.00112f
C248 adder_3_0/P4 CO 6.01e-19
C249 B1 adder_3_0/P2 6.78e-19
C250 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# -4.45e-20
C251 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# adder_3_0/P4 2.55e-19
C252 adder_3_0/G3 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 0.0333f
C253 adder_3_0/G2 A1 0.00324f
C254 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 4.82e-20
C255 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_3_0/P1 5.85e-19
C256 adder_2_0/G4 adder_3_0/G2 7.19e-19
C257 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# B3 4.93e-21
C258 adder_3_0/P1 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 0.0283f
C259 adder_3_0/P1 GND 0.175f
C260 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_3_0/P3 5.59e-20
C261 adder_3_0/P4 GND 0.492f
C262 adder_3_0/P1 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# 0.00281f
C263 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 0.00309f
C264 adder_3_0/P3 B2 0.00568f
C265 A2 A3 0.00214f
C266 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_3_0/P3 0.131f
C267 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.0026f
C268 adder_2_0/G4 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 4.89e-20
C269 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_3_0/sky130_fd_sc_hd__xor2_1_2/B -2.45e-19
C270 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X A3 5.54e-20
C271 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_117_297# adder_2_0/G4 3.36e-19
C272 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_3_0/P1 0.0152f
C273 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# B2 7.88e-20
C274 B4 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 5.38e-20
C275 adder_3_0/G3 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 3.99e-20
C276 VDD adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 5.68e-32
C277 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# VDD -5.68e-32
C278 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# B4 -3.44e-20
C279 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_47# adder_3_0/P3 -3.53e-19
C280 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 2.82e-21
C281 adder_3_0/P2 adder_3_0/G2 0.749f
C282 adder_3_0/P3 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# 1.03e-19
C283 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_3_0/P1 -9.58e-19
C284 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_3_0/P4 1.49e-19
C285 CO CI 0.0904f
C286 adder_3_0/G3 adder_2_0/sky130_fd_sc_hd__and4_1_0/X 4.68e-20
C287 adder_3_0/P1 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 0.00383f
C288 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# CI 0.0104f
C289 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_3_0/G2 0.00133f
C290 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# adder_3_0/G2 2.92e-19
C291 adder_2_0/sky130_fd_sc_hd__and4_1_0/X adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 6.99e-21
C292 adder_3_0/P2 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 0.00223f
C293 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_47# adder_3_0/sky130_fd_sc_hd__xor2_1_2/B -5.8e-19
C294 A1 B2 9.29e-19
C295 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# CI 2.49e-19
C296 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_2_0/G4 1.82e-19
C297 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B S3 -1.33e-20
C298 CO adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 6.62e-19
C299 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X CI 0.00101f
C300 B4 A4 1.95f
C301 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_117_297# S4 -3.24e-19
C302 adder_2_0/G4 B2 0.00161f
C303 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_3_0/sky130_fd_sc_hd__xor2_1_3/B -8.72e-21
C304 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_2_0/G4 1.36e-19
C305 GND CI 1.48f
C306 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# CI 4.51e-20
C307 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# adder_3_0/P1 1.85e-21
C308 VDD adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 1.34e-19
C309 B4 VDD 0.138f
C310 adder_3_0/P4 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 4.86e-19
C311 A3 adder_2_0/sky130_fd_sc_hd__and4_1_0/X 3.53e-20
C312 B4 B3 8.66e-19
C313 adder_3_0/G3 S1 6.53e-19
C314 adder_3_0/P3 A2 2.27e-19
C315 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X adder_3_0/P3 0.0225f
C316 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# CI 4.64e-20
C317 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# VDD -0.00753f
C318 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B S2 0.0038f
C319 S1 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.0236f
C320 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_47# S3 7.3e-19
C321 adder_3_0/G3 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 0.0407f
C322 adder_3_0/G3 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# -5.99e-22
C323 CO adder_2_0/sky130_fd_sc_hd__and4_1_0/a_303_47# 5.64e-19
C324 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# A2 1.08e-19
C325 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 0.00475f
C326 adder_2_0/G4 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# 5.98e-20
C327 adder_3_0/G2 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 9.85e-20
C328 adder_3_0/G3 adder_3_0/G1 0.0163f
C329 B1 A4 3.49e-19
C330 adder_3_0/P2 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 1.21e-19
C331 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_3_0/P3 0.00801f
C332 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# CI 0.00503f
C333 adder_3_0/G1 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B -6.76e-19
C334 B1 VDD 0.244f
C335 adder_3_0/P2 B2 0.0325f
C336 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_3_0/P2 0.0337f
C337 B1 B3 5.26e-19
C338 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# adder_3_0/P1 0.00658f
C339 S1 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_117_297# -4.4e-19
C340 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# CI 2.82e-19
C341 adder_3_0/P4 adder_3_0/P1 0.0308f
C342 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_384_47# adder_3_0/G1 1.56e-20
C343 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_3_0/G2 0.00912f
C344 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# VDD 0.00637f
C345 adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# B4 5.56e-19
C346 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# B2 0.00715f
C347 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_3_0/G2 1.11e-21
C348 A2 A1 0.00288f
C349 adder_3_0/P3 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 0.00835f
C350 A3 adder_3_0/G1 1.32e-19
C351 adder_2_0/G4 A2 1.33e-19
C352 adder_3_0/G3 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 0.00552f
C353 CI adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 0.00313f
C354 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 6.84e-21
C355 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X adder_2_0/G4 0.0203f
C356 adder_3_0/P2 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# -8.74e-21
C357 adder_3_0/P3 adder_2_0/sky130_fd_sc_hd__and4_1_0/X 5.85e-19
C358 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_384_47# adder_3_0/P1 5.17e-19
C359 S1 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 3.79e-19
C360 adder_3_0/G2 A4 1.16e-19
C361 adder_2_0/G4 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_47# 6.97e-19
C362 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_2_0/G4 1.01e-20
C363 VDD adder_3_0/G2 0.293f
C364 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 6.98e-20
C365 adder_3_0/G2 B3 1.49e-19
C366 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# B2 8.1e-20
C367 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# A4 3.72e-20
C368 adder_3_0/P3 S1 0.1f
C369 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# CI 0.0137f
C370 adder_3_0/P1 CI 0.154f
C371 adder_3_0/P4 CI 0.0664f
C372 adder_3_0/P2 A2 0.00581f
C373 VDD adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 3.32e-19
C374 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# B3 4.89e-20
C375 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X adder_3_0/P2 0.0208f
C376 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 8.63e-21
C377 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# adder_2_0/G4 1.75e-19
C378 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_109_47# adder_3_0/P3 4.98e-19
C379 CO adder_3_0/G3 4.09e-20
C380 adder_3_0/P3 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 0.024f
C381 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# adder_3_0/G3 3.83e-19
C382 adder_3_0/P3 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 3.07e-20
C383 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# B2 0.0195f
C384 S4 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.0035f
C385 CO adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.477f
C386 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 7.13e-21
C387 adder_3_0/P4 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 0.00212f
C388 adder_3_0/G3 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 0.00131f
C389 adder_3_0/P3 adder_3_0/G1 8.5e-20
C390 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_117_297# adder_3_0/G2 4.07e-19
C391 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_117_297# adder_3_0/P4 0.00227f
C392 adder_2_0/G4 adder_2_0/sky130_fd_sc_hd__and4_1_0/X 1.36e-19
C393 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_2_0/sky130_fd_sc_hd__and4_1_0/X 6.46e-21
C394 adder_3_0/G3 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 0.00133f
C395 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_3_0/sky130_fd_sc_hd__xor2_1_2/B -0.00531f
C396 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_3_0/P2 -8.11e-19
C397 adder_3_0/G3 GND 1.22f
C398 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_384_47# CI 2.66e-19
C399 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 1.8e-19
C400 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B GND -0.00596f
C401 CO A3 0.00124f
C402 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# adder_3_0/G1 0.0212f
C403 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# A3 2.34e-21
C404 adder_2_0/sky130_fd_sc_hd__and4_1_0/X S2 1.66e-20
C405 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# S3 -7.21e-19
C406 CO adder_2_0/sky130_fd_sc_hd__and4_1_0/a_197_47# 4.68e-19
C407 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# A4 3.72e-20
C408 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_47# S2 9.42e-19
C409 CO adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_117_297# 0.00216f
C410 adder_3_0/P3 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# -0.00186f
C411 adder_3_0/G3 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.00129f
C412 B4 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 0.0072f
C413 A4 B2 8.41e-19
C414 S1 S3 0.0279f
C415 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# VDD 2.99e-19
C416 adder_3_0/P2 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 4.11e-19
C417 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# B3 4.65e-20
C418 adder_2_0/G4 S1 2.86e-20
C419 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B S1 0.0151f
C420 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# adder_3_0/G2 2.56e-19
C421 adder_3_0/P3 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 0.0105f
C422 VDD B2 0.176f
C423 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B VDD -0.0577f
C424 A1 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 2.52e-21
C425 A3 GND 0.00693f
C426 B2 B3 0.00119f
C427 A2 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 9.74e-19
C428 adder_2_0/G4 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 0.0203f
C429 adder_3_0/P2 adder_2_0/sky130_fd_sc_hd__and4_1_0/X -2.14e-20
C430 adder_2_0/G4 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 0.00895f
C431 B1 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0.00727f
C432 A1 adder_3_0/G1 0.0955f
C433 B1 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# 0.00429f
C434 S1 S2 1.02f
C435 adder_3_0/G3 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 0.00395f
C436 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# A3 1e-19
C437 adder_2_0/G4 adder_3_0/G1 3.67e-20
C438 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_3_0/sky130_fd_sc_hd__xor2_1_2/B -0.00268f
C439 A2 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 1.78e-19
C440 CO adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 7.73e-19
C441 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 3.66e-20
C442 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 3.35e-21
C443 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# B3 0.00199f
C444 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_117_297# B2 0.00385f
C445 adder_3_0/G3 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 4.76e-20
C446 adder_3_0/P2 S1 0.234f
C447 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# S3 0.00612f
C448 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# GND 6.56e-19
C449 adder_3_0/G3 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 1.39e-19
C450 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# adder_3_0/sky130_fd_sc_hd__xor2_1_2/B -0.00349f
C451 adder_2_0/G4 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 1.03e-19
C452 S4 adder_3_0/P3 -8.8e-19
C453 CO adder_3_0/P3 0.0888f
C454 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# adder_3_0/P3 1.34e-19
C455 adder_3_0/P2 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 0.0193f
C456 B1 B4 2.5e-19
C457 A2 A4 4.9e-19
C458 adder_3_0/P3 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 1.7e-19
C459 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# S2 2.81e-19
C460 adder_3_0/P2 adder_3_0/G1 0.268f
C461 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 6.41e-20
C462 adder_3_0/G2 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 1.95e-19
C463 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# adder_3_0/G2 7.19e-20
C464 adder_3_0/P3 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 0.00384f
C465 A2 VDD 0.227f
C466 A2 B3 7.94e-19
C467 adder_3_0/P3 GND 0.136f
C468 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X VDD 0.00224f
C469 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 1.5e-20
C470 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_47# adder_3_0/G1 6.94e-19
C471 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X B3 1.6e-20
C472 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_3_0/G1 0.017f
C473 adder_3_0/G3 adder_3_0/P1 0.197f
C474 adder_3_0/P4 adder_3_0/G3 0.00126f
C475 adder_3_0/P2 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_384_47# 4.8e-19
C476 adder_3_0/P3 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 5.23e-19
C477 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# adder_3_0/sky130_fd_sc_hd__xor2_1_2/B -0.00512f
C478 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# GND 1.84e-20
C479 adder_3_0/P1 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.103f
C480 adder_3_0/P4 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 4.82e-19
C481 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# 6.41e-20
C482 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# VDD 3.54e-19
C483 S4 S3 0.442f
C484 adder_3_0/P2 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 0.00242f
C485 B1 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 8.1e-20
C486 CO S3 0.119f
C487 S4 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 0.00146f
C488 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# 1.09e-19
C489 CO adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 0.0228f
C490 CO adder_2_0/G4 1.56e-19
C491 B4 adder_3_0/G2 9.64e-20
C492 adder_3_0/G2 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 1.77e-21
C493 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 1.37e-21
C494 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# adder_2_0/G4 1.75e-19
C495 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_3_0/P3 1.78e-19
C496 A3 adder_3_0/P1 1.31e-19
C497 adder_3_0/P4 A3 1.54e-19
C498 adder_3_0/P3 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 5.91e-19
C499 adder_3_0/P1 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_197_47# 2.07e-19
C500 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X A1 2.97e-19
C501 adder_3_0/P4 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_117_297# 1.04e-19
C502 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# VDD 0.00235f
C503 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# adder_3_0/G2 3.05e-20
C504 A1 GND 0.00365f
C505 S4 S2 0.0289f
C506 CO S2 0.0426f
C507 S3 GND 0.0872f
C508 B4 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 3.05e-20
C509 adder_2_0/G4 GND 0.132f
C510 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B GND 0.00142f
C511 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_117_297# B4 0.00366f
C512 adder_2_0/sky130_fd_sc_hd__and4_1_0/X VDD -0.0032f
C513 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# adder_3_0/P3 0.00176f
C514 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# A1 -6.08e-19
C515 adder_2_0/sky130_fd_sc_hd__and4_1_0/X B3 1.55e-20
C516 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_145_75# adder_3_0/G2 8.25e-19
C517 adder_3_0/P3 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 1.36e-19
C518 B1 adder_3_0/G2 0.00409f
C519 S2 GND 0.089f
C520 adder_3_0/G3 CI 0.164f
C521 CO adder_3_0/P2 0.108f
C522 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_145_75# VDD 8.07e-19
C523 adder_3_0/P2 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_47# 0.00105f
C524 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# adder_3_0/P2 0.00114f
C525 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B CI -0.005f
C526 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_3_0/G2 0.00723f
C527 adder_3_0/P4 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 0.00101f
C528 adder_3_0/P2 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 0.00225f
C529 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_384_47# CI 1.5e-20
C530 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# A1 0.00131f
C531 S1 VDD -0.00144f
C532 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_2_0/G4 1.23e-20
C533 adder_3_0/P2 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 0.00437f
C534 adder_3_0/P2 GND 0.0707f
C535 adder_3_0/P2 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# 0.00724f
C536 B4 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 3.05e-20
C537 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# A4 -2.86e-19
C538 A3 CI 0.0954f
C539 VDD adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 0.00147f
C540 adder_3_0/P3 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# 1.5e-20
C541 B4 B2 4.83e-19
C542 VDD adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# -9.12e-19
C543 A4 adder_3_0/G1 7.97e-20
C544 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 2.14e-20
C545 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# -8.36e-21
C546 adder_3_0/P3 adder_3_0/P1 0.649f
C547 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_47# CI 9.49e-19
C548 adder_3_0/P4 adder_3_0/P3 0.232f
C549 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# GND 4.5e-19
C550 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# S2 0.00567f
C551 adder_3_0/P2 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 2.17e-19
C552 VDD adder_3_0/G1 0.694f
C553 adder_3_0/G1 B3 1.01e-19
C554 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# -0.00611f
C555 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# adder_3_0/P1 -6e-21
C556 A2 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# 5.47e-19
C557 A2 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0.00352f
C558 B1 B2 0.00145f
C559 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# adder_3_0/G2 1.78e-20
C560 adder_3_0/P2 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# -1.88e-20
C561 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_384_47# adder_3_0/G2 7.32e-20
C562 adder_3_0/P1 A1 0.00472f
C563 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# GND 1.04e-19
C564 adder_3_0/P4 S3 0.0135f
C565 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# adder_3_0/P2 0.00898f
C566 adder_2_0/G4 adder_3_0/P1 0.03f
C567 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_3_0/P1 -6.47e-19
C568 adder_3_0/P4 adder_2_0/G4 1.29f
C569 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# S1 -1.39e-20
C570 adder_3_0/P4 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 0.0108f
C571 adder_3_0/P3 CI 0.132f
C572 B4 A2 3.27e-19
C573 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# GND -2.23e-19
C574 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 9.82e-21
C575 adder_3_0/P4 S2 9.76e-19
C576 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# GND -2.36e-19
C577 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 1.53e-19
C578 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_3_0/G2 0.0173f
C579 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# adder_3_0/P3 3.13e-19
C580 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# CI 2.96e-20
C581 adder_3_0/G2 B2 0.089f
C582 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_3_0/G2 0.0309f
C583 S4 VDD -2.22e-19
C584 CO VDD 0.114f
C585 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# VDD 0.00215f
C586 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# B3 9.41e-19
C587 adder_3_0/P2 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# 0.00132f
C588 adder_3_0/P4 adder_3_0/P2 0.0172f
C589 adder_3_0/P2 adder_3_0/P1 1.17f
C590 B1 A2 0.403f
C591 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# VDD 6.69e-20
C592 A4 GND 0.00516f
C593 adder_3_0/P3 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_303_47# 4e-19
C594 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_47# adder_3_0/P1 0.00105f
C595 VDD adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 0.0342f
C596 A1 CI 1.72e-19
C597 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# adder_3_0/P1 3.68e-21
C598 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_3_0/P1 7.78e-20
C599 adder_3_0/G3 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.00104f
C600 adder_3_0/P4 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 2.19e-20
C601 VDD GND 1.2f
C602 B3 GND 0.00596f
C603 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B CI 1.31e-19
C604 adder_2_0/G4 CI 0.0329f
C605 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# A4 6.49e-20
C606 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# VDD -4.41e-19
C607 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# B3 7.98e-20
C608 adder_3_0/G3 A3 0.0807f
C609 S2 CI 0.00387f
C610 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_117_297# adder_2_0/G4 3.67e-19
C611 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# adder_3_0/G1 3.22e-19
C612 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# adder_3_0/G1 4.07e-19
C613 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# B2 6.16e-19
C614 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# VDD 4.68e-19
C615 A2 adder_3_0/G2 0.084f
C616 VDD adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 0.00221f
C617 adder_3_0/P1 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 5.66e-20
C618 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X adder_3_0/G2 1.74e-19
C619 adder_3_0/P4 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 4.73e-19
C620 adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# GND 3.16e-20
C621 S1 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# -1.76e-19
C622 adder_3_0/P2 CI 0.0316f
C623 CO adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# 4.34e-19
C624 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# CI 0.0052f
C625 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# S1 -2.34e-19
C626 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 9.58e-21
C627 B4 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 0.0208f
C628 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# GND -5.95e-20
C629 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_3_0/P1 1.38e-19
C630 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 8.48e-19
C631 adder_3_0/P4 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 7.7e-20
C632 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 2.84e-32
C633 adder_3_0/P4 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 5.92e-20
C634 B4 adder_3_0/G1 6.45e-20
C635 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 2.99e-20
C636 adder_3_0/G3 adder_3_0/P3 0.318f
C637 adder_3_0/P2 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_303_47# 1.69e-19
C638 adder_3_0/P3 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.00276f
C639 B1 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 3.97e-19
C640 adder_3_0/P1 A4 8.78e-20
C641 adder_3_0/P4 A4 0.00541f
C642 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# GND -5.69e-20
C643 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# A2 0.0155f
C644 B1 adder_3_0/G1 0.087f
C645 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# CI 2.83e-19
C646 VDD adder_3_0/P1 0.332f
C647 adder_3_0/P4 VDD 0.896f
C648 adder_3_0/P1 B3 1.06e-19
C649 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 2.6e-21
C650 A2 B2 0.77f
C651 adder_3_0/P4 B3 1.46e-19
C652 CO adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0.00661f
C653 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_3_0/G1 0.0239f
C654 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X B2 1.92e-20
C655 adder_3_0/P3 A3 0.002f
C656 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 1.11e-19
C657 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_145_75# adder_3_0/G2 5.09e-21
C658 adder_3_0/P3 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_197_47# 4.99e-19
C659 adder_3_0/P3 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_47# 9.41e-19
C660 adder_3_0/P3 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_117_297# 1.69e-19
C661 adder_2_0/sky130_fd_sc_hd__and4_1_0/X adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 7.41e-22
C662 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# CI 4.53e-20
C663 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# CI 0.0185f
C664 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# A3 5.96e-20
C665 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# -9.51e-19
C666 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# 4.7e-20
C667 adder_3_0/G3 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 0.0127f
C668 adder_3_0/G3 adder_2_0/G4 0.217f
C669 adder_3_0/P1 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_117_297# 3.02e-21
C670 S3 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.0023f
C671 adder_3_0/G2 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 0.0356f
C672 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_3_0/sky130_fd_sc_hd__xor2_1_2/B -0.0029f
C673 adder_2_0/G4 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 8.62e-20
C674 adder_3_0/P4 adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 4.95e-20
C675 adder_3_0/P3 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 2.95e-20
C676 adder_3_0/G2 adder_3_0/G1 0.872f
C677 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# B2 5.71e-20
C678 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 1.39e-20
C679 A4 CI 0.0346f
C680 A3 A1 5.77e-19
C681 CO adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# 8.7e-19
C682 S2 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0.118f
C683 CO adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 1.62e-20
C684 adder_3_0/P3 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_47# 1.14e-19
C685 VDD CI 1.6f
C686 adder_2_0/G4 A3 2.73e-19
C687 B3 CI 0.208f
C688 adder_3_0/P4 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# -2.02e-20
C689 B4 GND 0.00678f
C690 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# GND 4.59e-19
C691 adder_3_0/P4 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 0.0105f
C692 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_2_0/sky130_fd_sc_hd__and4_1_0/X 7.03e-19
C693 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_384_47# adder_3_0/G2 4.16e-19
C694 adder_3_0/P4 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_117_297# 4.5e-19
C695 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X A2 2.61e-19
C696 adder_3_0/G3 adder_3_0/P2 0.771f
C697 adder_3_0/P2 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B -0.0409f
C698 B4 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 5.38e-20
C699 adder_3_0/G3 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_47# 0.00103f
C700 adder_3_0/G3 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 1.82e-20
C701 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_3_0/sky130_fd_sc_hd__xor2_1_2/B -0.00197f
C702 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B S1 0.00968f
C703 B1 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 2.31e-20
C704 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# S3 0.00559f
C705 adder_3_0/P1 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# 0.00143f
C706 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 9.34e-21
C707 adder_3_0/P4 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# 1.73e-19
C708 B1 GND 0.00716f
C709 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 4.59e-19
C710 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# -0.00152f
C711 adder_2_0/G4 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 3.23e-20
C712 adder_3_0/P2 A3 0.0346f
C713 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_47# S3 9.42e-19
C714 B2 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 2.07e-20
C715 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 5.75e-20
C716 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# GND 9.07e-20
C717 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# adder_3_0/G1 3.92e-20
C718 A3 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 9.09e-19
C719 B1 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 0.022f
C720 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# S2 0.00273f
C721 B2 adder_3_0/G1 2.02e-19
C722 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_3_0/G1 0.0407f
C723 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# -1.77e-19
C724 adder_3_0/P3 S3 0.0899f
C725 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# CI 0.00281f
C726 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_3_0/P3 -0.00685f
C727 adder_3_0/P3 adder_2_0/G4 1.15f
C728 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_47# adder_3_0/G2 6.94e-19
C729 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_117_297# adder_3_0/P1 3.41e-19
C730 adder_3_0/G3 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0.0177f
C731 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# adder_3_0/P1 5.1e-19
C732 adder_3_0/P1 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0.00383f
C733 adder_3_0/G3 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_145_75# 8.23e-19
C734 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X adder_2_0/sky130_fd_sc_hd__and4_1_0/X -0.0153f
C735 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# A1 0.0155f
C736 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_384_47# 7.89e-20
C737 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 4.77e-19
C738 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# adder_3_0/G2 0.0146f
C739 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 0.00238f
C740 B1 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 3.89e-20
C741 adder_3_0/P2 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# -4.84e-19
C742 adder_3_0/P3 S2 0.238f
C743 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# -3.51e-21
C744 adder_3_0/P4 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 0.011f
C745 adder_3_0/G2 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 0.0275f
C746 CO adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 4.8e-20
C747 adder_3_0/G2 GND 0.287f
C748 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 1.13e-19
C749 adder_3_0/G2 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# 0.0051f
C750 adder_3_0/G3 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 4.15e-19
C751 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 2.85e-19
C752 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# adder_3_0/G3 0.00202f
C753 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# CI 0.0208f
C754 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X S1 6.31e-20
C755 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# adder_3_0/G2 0.00105f
C756 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# GND 3.52e-21
C757 adder_3_0/P2 adder_3_0/P3 0.405f
C758 B4 adder_3_0/P1 4.85e-20
C759 adder_3_0/P1 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 2.37e-21
C760 A2 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 1.47e-20
C761 adder_3_0/P4 B4 0.0321f
C762 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B S3 0.045f
C763 adder_2_0/G4 S3 2.78e-20
C764 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_3_0/P3 5.63e-21
C765 A3 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 5.49e-19
C766 adder_3_0/P3 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 1.27e-21
C767 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B adder_2_0/G4 0.00256f
C768 A2 adder_3_0/G1 3.33e-19
C769 adder_3_0/P4 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 5.12e-19
C770 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# S1 5.99e-19
C771 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# A3 -7.46e-20
C772 adder_3_0/G3 A4 1.67e-19
C773 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X adder_3_0/G1 3.53e-20
C774 adder_3_0/G2 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 0.0185f
C775 adder_3_0/G3 VDD 0.253f
C776 S2 S3 0.717f
C777 adder_3_0/G3 B3 0.0363f
C778 adder_2_0/G4 S2 2.28e-20
C779 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B S2 0.0283f
C780 VDD adder_3_0/sky130_fd_sc_hd__xor2_1_2/B -0.019f
C781 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B CO 0.0577f
C782 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# 0.00254f
C783 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_145_75# adder_3_0/P1 6.85e-19
C784 B1 adder_3_0/P1 0.0278f
C785 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# S1 9.19e-19
C786 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# adder_3_0/G2 0.00591f
C787 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# GND 1.84e-20
C788 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# adder_3_0/P1 0.00259f
C789 adder_3_0/P2 A1 3.75e-19
C790 A3 A4 0.00106f
C791 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 0 0.00137f
C792 adder_1_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 0 0.255f
C793 A2 0 0.553f
C794 B2 0 0.632f
C795 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 0 0.00137f
C796 adder_1_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 0 0.255f
C797 A1 0 0.469f
C798 B1 0 0.496f
C799 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0 0.00137f
C800 adder_1_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 0 0.255f
C801 B4 0 1.05f
C802 A4 0 0.714f
C803 adder_1_0/sky130_fd_sc_hd__and2_1_3/a_59_75# 0 0.177f
C804 B3 0 0.683f
C805 A3 0 0.729f
C806 adder_1_0/sky130_fd_sc_hd__and2_1_2/a_59_75# 0 0.177f
C807 adder_1_0/sky130_fd_sc_hd__and2_1_1/a_59_75# 0 0.177f
C808 adder_1_0/sky130_fd_sc_hd__and2_1_0/a_59_75# 0 0.177f
C809 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 0 0.00137f
C810 adder_1_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 0 0.255f
C811 S3 0 0.233f
C812 adder_3_0/P3 0 1.49f
C813 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_285_297# 0 0.00137f
C814 adder_3_0/sky130_fd_sc_hd__xor2_1_2/a_35_297# 0 0.255f
C815 GND 0 9.62f
C816 S2 0 0.212f
C817 adder_3_0/P2 0 1.26f
C818 adder_3_0/sky130_fd_sc_hd__xor2_1_1/B 0 0.486f
C819 VDD 0 17.4f
C820 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_285_297# 0 0.00137f
C821 adder_3_0/sky130_fd_sc_hd__xor2_1_1/a_35_297# 0 0.255f
C822 S1 0 0.353f
C823 adder_3_0/P1 0 1.11f
C824 CI 0 2.13f
C825 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_285_297# 0 0.00137f
C826 adder_3_0/sky130_fd_sc_hd__xor2_1_0/a_35_297# 0 0.255f
C827 adder_3_0/sky130_fd_sc_hd__xor2_1_3/B 0 0.336f
C828 adder_3_0/sky130_fd_sc_hd__xor2_1_2/B 0 1.53f
C829 adder_3_0/G3 0 0.718f
C830 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 0 0.0348f
C831 adder_3_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0 0.147f
C832 adder_3_0/G2 0 0.642f
C833 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 0 0.0348f
C834 adder_3_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 0 0.147f
C835 adder_3_0/G1 0 0.527f
C836 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# 0 0.0348f
C837 adder_3_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 0 0.147f
C838 S4 0 0.344f
C839 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_285_297# 0 0.00137f
C840 adder_3_0/sky130_fd_sc_hd__xor2_1_3/a_35_297# 0 0.255f
C841 adder_2_0/sky130_fd_sc_hd__and4_1_0/X 0 0.154f
C842 adder_3_0/P4 0 1.62f
C843 adder_2_0/sky130_fd_sc_hd__and4_1_0/a_27_47# 0 0.175f
C844 CO 0 0.959f
C845 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_299_297# 0 0.0348f
C846 adder_2_0/sky130_fd_sc_hd__a21o_1_3/a_81_21# 0 0.147f
C847 adder_2_0/sky130_fd_sc_hd__a21o_1_2/X 0 0.168f
C848 adder_2_0/sky130_fd_sc_hd__a21o_1_1/X 0 0.129f
C849 adder_2_0/G4 0 0.596f
C850 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_299_297# 0 0.0348f
C851 adder_2_0/sky130_fd_sc_hd__a21o_1_2/a_81_21# 0 0.147f
C852 adder_2_0/sky130_fd_sc_hd__a21o_1_0/X 0 0.223f
C853 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_299_297# 0 0.0348f
C854 adder_2_0/sky130_fd_sc_hd__a21o_1_1/a_81_21# 0 0.147f
C855 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_299_297# 0 0.0348f
C856 adder_2_0/sky130_fd_sc_hd__a21o_1_0/a_81_21# 0 0.147f
.ends

.GLOBAL GND

.end

