magic
tech sky130A
magscale 1 2
timestamp 1701618932
<< metal1 >>
rect 3290 1445 3370 1455
rect 3290 1430 3300 1445
rect 15 1400 3300 1430
rect 3290 1385 3300 1400
rect 3360 1385 3370 1445
rect 3290 1375 3370 1385
rect 4630 1360 4710 1370
rect 4630 1345 4640 1360
rect 15 1315 4640 1345
rect 4630 1300 4640 1315
rect 4700 1300 4710 1360
rect 4630 1290 4710 1300
rect 4065 1275 4145 1285
rect 4065 1260 4075 1275
rect 15 1230 4075 1260
rect 4065 1215 4075 1230
rect 4135 1215 4145 1275
rect 4065 1205 4145 1215
rect 3600 1190 3680 1200
rect 3600 1175 3610 1190
rect 15 1145 3610 1175
rect 3600 1130 3610 1145
rect 3670 1130 3680 1190
rect 3600 1120 3680 1130
rect 2785 1105 2865 1115
rect 2785 1090 2795 1105
rect 15 1060 2795 1090
rect 2785 1045 2795 1060
rect 2855 1045 2865 1105
rect 2785 1035 2865 1045
rect 1910 1020 1990 1030
rect 1910 1005 1920 1020
rect 15 975 1920 1005
rect 1910 960 1920 975
rect 1980 960 1990 1020
rect 1910 950 1990 960
rect 1350 935 1425 945
rect 1350 920 1360 935
rect 15 890 1360 920
rect 1350 875 1360 890
rect 1415 875 1425 935
rect 1350 865 1425 875
rect 635 850 715 860
rect 635 835 645 850
rect 15 805 645 835
rect 635 790 645 805
rect 705 790 715 850
rect 635 780 715 790
rect 70 765 150 775
rect 70 750 80 765
rect 15 720 80 750
rect 70 705 80 720
rect 140 705 150 765
rect 70 695 150 705
rect 360 510 440 520
rect 360 450 370 510
rect 430 450 440 510
rect 360 440 440 450
rect 1640 515 1720 525
rect 1640 455 1650 515
rect 1710 455 1720 515
rect 1640 445 1720 455
rect 2390 500 2470 510
rect 1110 435 1190 445
rect 1110 375 1120 435
rect 1180 375 1190 435
rect 2390 440 2400 500
rect 2460 440 2470 500
rect 2390 430 2470 440
rect 3080 505 3160 515
rect 3080 445 3090 505
rect 3150 445 3160 505
rect 3080 435 3160 445
rect 4360 510 4435 520
rect 4360 450 4370 510
rect 4425 450 4435 510
rect 4360 440 4435 450
rect 5110 495 5190 505
rect 3830 430 3910 440
rect 1110 365 1190 375
rect 3830 370 3840 430
rect 3900 370 3910 430
rect 5110 435 5120 495
rect 5180 435 5190 495
rect 5110 425 5190 435
rect 3830 360 3910 370
rect 360 -15 440 -5
rect 360 -30 370 -15
rect 50 -60 370 -30
rect 360 -75 370 -60
rect 430 -75 440 -15
rect 360 -85 440 -75
rect 860 -15 940 -5
rect 860 -75 870 -15
rect 930 -30 940 -15
rect 3080 -15 3160 -5
rect 3080 -30 3090 -15
rect 930 -60 3090 -30
rect 930 -75 940 -60
rect 860 -85 940 -75
rect 3080 -75 3090 -60
rect 3150 -75 3160 -15
rect 3080 -85 3160 -75
rect 220 -100 300 -90
rect 220 -115 230 -100
rect 120 -145 230 -115
rect 220 -160 230 -145
rect 290 -115 300 -100
rect 1640 -100 1720 -90
rect 1640 -115 1650 -100
rect 290 -145 1650 -115
rect 290 -160 300 -145
rect 220 -170 300 -160
rect 1640 -160 1650 -145
rect 1710 -160 1720 -100
rect 1640 -170 1720 -160
rect 475 -185 555 -175
rect 475 -245 485 -185
rect 545 -200 555 -185
rect 2390 -185 2470 -175
rect 2390 -200 2400 -185
rect 545 -230 2400 -200
rect 545 -245 555 -230
rect 475 -255 555 -245
rect 2390 -245 2400 -230
rect 2460 -245 2470 -185
rect 2390 -255 2470 -245
rect 1110 -295 1190 -285
rect 1110 -310 1120 -295
rect 585 -340 1120 -310
rect 1110 -355 1120 -340
rect 1180 -310 1190 -295
rect 2470 -295 2550 -285
rect 2470 -310 2480 -295
rect 1180 -340 2480 -310
rect 1180 -355 1190 -340
rect 1110 -365 1190 -355
rect 2470 -355 2480 -340
rect 2540 -355 2550 -295
rect 2470 -365 2550 -355
rect 1115 -405 1195 -395
rect 1115 -465 1125 -405
rect 1185 -420 1195 -405
rect 3830 -405 3910 -395
rect 3830 -420 3840 -405
rect 1185 -450 3840 -420
rect 1185 -465 1195 -450
rect 1115 -475 1195 -465
rect 3830 -465 3840 -450
rect 3900 -465 3910 -405
rect 3830 -475 3910 -465
rect 1500 -490 1580 -480
rect 1500 -550 1510 -490
rect 1570 -505 1580 -490
rect 4360 -490 4440 -480
rect 4360 -505 4370 -490
rect 1570 -535 4370 -505
rect 1570 -550 1580 -535
rect 1500 -560 1580 -550
rect 4360 -550 4370 -535
rect 4430 -550 4440 -490
rect 4360 -560 4440 -550
rect 1760 -575 1840 -565
rect 1760 -630 1770 -575
rect 1830 -590 1840 -575
rect 5110 -575 5190 -565
rect 5110 -590 5120 -575
rect 1830 -620 5120 -590
rect 1830 -630 1840 -620
rect 1760 -640 1840 -630
rect 5110 -635 5120 -620
rect 5180 -635 5190 -575
rect 5110 -645 5190 -635
rect 3295 -1005 3375 -995
rect 1115 -1080 1195 -1005
rect 3295 -1065 3305 -1005
rect 3365 -1065 3375 -1005
rect 3295 -1075 3375 -1065
rect 1115 -1085 1120 -1080
rect 1140 -1085 1195 -1080
rect 345 -1360 425 -1350
rect 345 -1420 355 -1360
rect 415 -1375 425 -1360
rect 3295 -1360 3375 -1350
rect 3295 -1375 3305 -1360
rect 415 -1405 3305 -1375
rect 415 -1420 425 -1405
rect 345 -1430 425 -1420
rect 3295 -1420 3305 -1405
rect 3365 -1420 3375 -1360
rect 3295 -1430 3375 -1420
rect 1745 -1599 1825 -1589
rect 1745 -1659 1755 -1599
rect 1815 -1614 1825 -1599
rect 1900 -1599 1980 -1589
rect 1900 -1614 1910 -1599
rect 1815 -1644 1910 -1614
rect 1815 -1659 1825 -1644
rect 1745 -1669 1825 -1659
rect 1900 -1659 1910 -1644
rect 1970 -1659 1980 -1599
rect 1900 -1669 1980 -1659
rect 3265 -2155 3345 -2130
rect 3265 -2185 5590 -2155
rect 3265 -2210 3345 -2185
rect 3990 -2225 4070 -2215
rect 3990 -2285 4000 -2225
rect 4060 -2240 4070 -2225
rect 4060 -2270 5590 -2240
rect 4060 -2285 4070 -2270
rect 3990 -2295 4070 -2285
rect 4720 -2310 4800 -2300
rect 4720 -2370 4730 -2310
rect 4790 -2325 4800 -2310
rect 4790 -2355 5590 -2325
rect 4790 -2370 4800 -2355
rect 4720 -2380 4800 -2370
rect 5450 -2395 5530 -2385
rect 5450 -2455 5460 -2395
rect 5520 -2410 5530 -2395
rect 5520 -2440 5590 -2410
rect 5520 -2455 5530 -2440
rect 5450 -2465 5530 -2455
rect 1930 -2650 2010 -2640
rect 1930 -2710 1940 -2650
rect 2000 -2665 2010 -2650
rect 2000 -2695 5590 -2665
rect 2000 -2710 2010 -2695
rect 1930 -2720 2010 -2710
<< via1 >>
rect 3300 1385 3360 1445
rect 4640 1300 4700 1360
rect 4075 1215 4135 1275
rect 3610 1130 3670 1190
rect 2795 1045 2855 1105
rect 1920 960 1980 1020
rect 1360 875 1415 935
rect 645 790 705 850
rect 80 705 140 765
rect 370 450 430 510
rect 1650 455 1710 515
rect 1120 375 1180 435
rect 2400 440 2460 500
rect 3090 445 3150 505
rect 4370 450 4425 510
rect 3840 370 3900 430
rect 5120 435 5180 495
rect 370 -75 430 -15
rect 870 -75 930 -15
rect 3090 -75 3150 -15
rect 230 -160 290 -100
rect 1650 -160 1710 -100
rect 485 -245 545 -185
rect 2400 -245 2460 -185
rect 1120 -355 1180 -295
rect 2480 -355 2540 -295
rect 1125 -465 1185 -405
rect 3840 -465 3900 -405
rect 1510 -550 1570 -490
rect 4370 -550 4430 -490
rect 1770 -630 1830 -575
rect 5120 -635 5180 -575
rect 3305 -1065 3365 -1005
rect 355 -1420 415 -1360
rect 3305 -1420 3365 -1360
rect 1755 -1659 1815 -1599
rect 1910 -1659 1970 -1599
rect 4000 -2285 4060 -2225
rect 4730 -2370 4790 -2310
rect 5460 -2455 5520 -2395
rect 1940 -2710 2000 -2650
<< metal2 >>
rect 3290 1445 3370 1455
rect 3290 1385 3300 1445
rect 3360 1385 3370 1445
rect 3290 1375 3370 1385
rect 2785 1105 2865 1115
rect 2785 1045 2795 1105
rect 2855 1045 2865 1105
rect 2785 1035 2865 1045
rect 1910 1020 1990 1030
rect 1910 960 1920 1020
rect 1980 960 1990 1020
rect 1910 950 1990 960
rect 1350 935 1425 945
rect 1350 875 1360 935
rect 1415 875 1425 935
rect 1350 865 1425 875
rect 635 850 715 860
rect 635 790 645 850
rect 705 790 715 850
rect 635 780 715 790
rect 70 765 150 775
rect 70 705 80 765
rect 140 705 150 765
rect 70 695 150 705
rect 95 325 125 695
rect 360 510 440 520
rect 360 450 370 510
rect 430 450 440 510
rect 360 440 440 450
rect 385 -5 415 440
rect 660 325 690 780
rect 1110 435 1190 445
rect 1110 375 1120 435
rect 1180 375 1190 435
rect 1110 365 1190 375
rect 360 -15 440 -5
rect 120 -1804 150 -15
rect 360 -75 370 -15
rect 430 -75 440 -15
rect 360 -85 440 -75
rect 860 -15 940 -5
rect 860 -75 870 -15
rect 930 -75 940 -15
rect 860 -85 940 -75
rect 220 -100 300 -90
rect 220 -160 230 -100
rect 290 -160 300 -100
rect 220 -170 300 -160
rect 245 -1010 275 -170
rect 370 -1010 400 -85
rect 475 -185 555 -175
rect 475 -245 485 -185
rect 545 -245 555 -185
rect 475 -255 555 -245
rect 500 -1010 530 -255
rect 215 -1050 225 -1020
rect 550 -1050 560 -1020
rect 245 -1085 275 -1075
rect 370 -1085 400 -1075
rect 500 -1085 530 -1070
rect 345 -1360 425 -1350
rect 345 -1420 355 -1360
rect 415 -1420 425 -1360
rect 345 -1430 425 -1420
rect 370 -1800 400 -1430
rect 600 -1799 630 -285
rect 120 -1834 225 -1804
rect 560 -1829 630 -1799
rect 775 -1804 805 -100
rect 885 -1015 915 -85
rect 1135 -285 1165 365
rect 1375 325 1405 865
rect 1640 515 1720 525
rect 1640 455 1650 515
rect 1710 455 1720 515
rect 1640 445 1720 455
rect 1110 -295 1190 -285
rect 1110 -355 1120 -295
rect 1180 -355 1190 -295
rect 1110 -365 1190 -355
rect 1115 -405 1195 -395
rect 1115 -465 1125 -405
rect 1185 -465 1195 -405
rect 1115 -475 1195 -465
rect 1140 -1005 1170 -475
rect 885 -1085 915 -1060
rect 1115 -1085 1195 -1005
rect 1140 -1090 1170 -1085
rect 1245 -1804 1275 -180
rect 775 -1834 860 -1804
rect 1190 -1834 1275 -1804
rect 1400 -1804 1430 -15
rect 1665 -90 1695 445
rect 1935 325 1965 950
rect 2390 500 2470 510
rect 2390 440 2400 500
rect 2460 440 2470 500
rect 2390 430 2470 440
rect 1640 -100 1720 -90
rect 1640 -160 1650 -100
rect 1710 -160 1720 -100
rect 1640 -170 1720 -160
rect 2415 -175 2445 430
rect 2810 325 2840 1035
rect 3080 505 3160 515
rect 3080 445 3090 505
rect 3150 445 3160 505
rect 3080 435 3160 445
rect 3105 -5 3135 435
rect 3080 -15 3160 -5
rect 3080 -75 3090 -15
rect 3150 -75 3160 -15
rect 3080 -85 3160 -75
rect 2390 -185 2470 -175
rect 2390 -245 2400 -185
rect 2460 -245 2470 -185
rect 2390 -255 2470 -245
rect 2470 -295 2550 -285
rect 2470 -355 2480 -295
rect 2540 -355 2550 -295
rect 2470 -365 2550 -355
rect 1500 -490 1580 -480
rect 1500 -550 1510 -490
rect 1570 -550 1580 -490
rect 1500 -560 1580 -550
rect 1525 -1015 1555 -560
rect 1760 -575 1840 -565
rect 1760 -630 1770 -575
rect 1830 -630 1840 -575
rect 1760 -640 1840 -630
rect 1785 -1015 1815 -640
rect 1525 -1080 1555 -1060
rect 1785 -1080 1815 -1065
rect 1925 -1589 1955 -395
rect 1745 -1599 1825 -1589
rect 1745 -1659 1755 -1599
rect 1815 -1659 1825 -1599
rect 1745 -1669 1825 -1659
rect 1900 -1599 1980 -1589
rect 1900 -1659 1910 -1599
rect 1970 -1659 1980 -1599
rect 1900 -1669 1980 -1659
rect 1770 -1799 1800 -1669
rect 2150 -1794 2180 -480
rect 2405 -1799 2435 -480
rect 2490 -1045 2520 -365
rect 3315 -995 3345 1375
rect 4630 1360 4710 1370
rect 4630 1300 4640 1360
rect 4700 1300 4710 1360
rect 4630 1290 4710 1300
rect 4065 1275 4145 1285
rect 4065 1215 4075 1275
rect 4135 1215 4145 1275
rect 4065 1205 4145 1215
rect 3600 1190 3680 1200
rect 3600 1130 3610 1190
rect 3670 1130 3680 1190
rect 3600 1120 3680 1130
rect 3625 325 3655 1120
rect 3830 430 3910 440
rect 3830 370 3840 430
rect 3900 370 3910 430
rect 3830 360 3910 370
rect 3855 -395 3885 360
rect 4090 325 4120 1205
rect 4360 510 4435 520
rect 4360 450 4370 510
rect 4425 450 4435 510
rect 4360 440 4435 450
rect 3830 -405 3910 -395
rect 3830 -465 3840 -405
rect 3900 -465 3910 -405
rect 3830 -475 3910 -465
rect 4385 -480 4415 440
rect 4655 325 4685 1290
rect 5110 495 5190 505
rect 5110 435 5120 495
rect 5180 435 5190 495
rect 5110 425 5190 435
rect 4360 -490 4440 -480
rect 4360 -550 4370 -490
rect 4430 -550 4440 -490
rect 4360 -560 4440 -550
rect 5135 -565 5165 425
rect 5110 -575 5190 -565
rect 5110 -635 5120 -575
rect 5180 -635 5190 -575
rect 5110 -645 5190 -635
rect 3295 -1005 3375 -995
rect 2490 -1090 2520 -1060
rect 3295 -1065 3305 -1005
rect 3365 -1065 3375 -1005
rect 3295 -1075 3375 -1065
rect 3320 -1350 3350 -1075
rect 3295 -1360 3375 -1350
rect 3295 -1420 3305 -1360
rect 3365 -1420 3375 -1360
rect 3295 -1430 3375 -1420
rect 1400 -1834 1495 -1804
rect 1955 -2640 1985 -1830
rect 3290 -2130 3320 -1760
rect 3265 -2210 3345 -2130
rect 4015 -2215 4045 -1745
rect 3990 -2225 4070 -2215
rect 3990 -2285 4000 -2225
rect 4060 -2285 4070 -2225
rect 3990 -2295 4070 -2285
rect 4745 -2300 4775 -1755
rect 4720 -2310 4800 -2300
rect 4720 -2370 4730 -2310
rect 4790 -2370 4800 -2310
rect 4720 -2380 4800 -2370
rect 5475 -2385 5505 -1745
rect 5450 -2395 5530 -2385
rect 5450 -2455 5460 -2395
rect 5520 -2455 5530 -2395
rect 5450 -2465 5530 -2455
rect 1930 -2650 2010 -2640
rect 1930 -2710 1940 -2650
rect 2000 -2710 2010 -2650
rect 1930 -2720 2010 -2710
use adder_1  adder_1_0
timestamp 1700079872
transform 1 0 60 0 1 74
box -80 -50 5188 590
use adder_2  adder_2_0
timestamp 1700046346
transform 1 0 30 0 1 -1277
box -50 -40 3394 600
use adder_3  adder_3_0
timestamp 1699994886
transform 1 0 25 0 1 -2055
box -45 -580 5561 595
<< end >>
