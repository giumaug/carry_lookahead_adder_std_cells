magic
tech sky130A
magscale 1 2
timestamp 1695416290
<< nwell >>
rect 433 259 473 580
rect 1184 259 1204 580
rect 1207 259 1247 579
rect 1724 259 1754 580
rect 2465 259 2483 580
rect 3009 259 3033 580
rect 3742 259 3763 580
rect 4288 259 4316 580
<< locali >>
rect 412 525 444 559
rect 480 525 513 559
rect 1144 525 1180 559
rect 1215 525 1245 559
rect 1693 525 1724 559
rect 1760 525 1793 559
rect 2426 525 2454 559
rect 2490 525 2523 559
rect 2974 525 3005 559
rect 3040 525 3073 559
rect 3704 525 3740 559
rect 3775 525 3804 559
rect 4253 525 4285 559
rect 4320 525 4354 559
rect 340 420 375 454
rect 397 -20 444 15
rect 480 -20 515 15
rect 1147 -19 1174 15
rect 1210 -19 1246 15
rect 1686 -19 1725 15
rect 1760 -19 1795 15
rect 2427 -19 2460 15
rect 2495 -19 2523 15
rect 2966 -19 3005 15
rect 3040 -19 3071 15
rect 3706 -19 3740 15
rect 3775 -19 3802 15
rect 4247 -19 4285 15
rect 4320 -19 4355 15
<< viali >>
rect 79 525 113 559
rect 444 525 480 559
rect 1180 525 1215 559
rect 1724 525 1760 559
rect 2454 525 2490 559
rect 3005 525 3040 559
rect 3740 525 3775 559
rect 4285 525 4320 559
rect 325 381 359 415
rect 1605 381 1639 415
rect 2355 373 2389 407
rect 2885 381 2919 415
rect 4165 381 4199 415
rect 4915 373 4949 407
rect 1075 305 1109 339
rect 3635 305 3669 339
rect 32 213 66 247
rect 173 213 207 247
rect 593 213 627 247
rect 710 213 744 247
rect 1312 213 1346 247
rect 1453 213 1487 247
rect 1873 213 1907 247
rect 1990 213 2024 247
rect 2592 213 2626 247
rect 2733 213 2767 247
rect 3270 213 3304 247
rect 3405 213 3439 247
rect 3872 213 3906 247
rect 4013 213 4047 247
rect 4433 213 4467 247
rect 4550 213 4584 247
rect 444 -20 480 15
rect 1174 -19 1210 15
rect 1725 -19 1760 15
rect 2460 -19 2495 15
rect 3005 -19 3040 15
rect 3740 -19 3775 15
rect 4285 -19 4320 15
<< metal1 >>
rect 413 559 511 590
rect 413 525 444 559
rect 480 525 511 559
rect 413 494 511 525
rect 1145 559 1242 590
rect 1145 525 1180 559
rect 1215 525 1242 559
rect 1145 494 1242 525
rect 1693 559 1791 590
rect 1693 525 1724 559
rect 1760 525 1791 559
rect 1693 494 1791 525
rect 2425 559 2522 590
rect 2425 525 2454 559
rect 2490 525 2522 559
rect 2425 494 2522 525
rect 2972 559 3073 590
rect 2972 525 3005 559
rect 3040 525 3073 559
rect 2972 494 3073 525
rect 3706 559 3804 590
rect 3706 525 3740 559
rect 3775 525 3804 559
rect 3706 494 3804 525
rect 4253 559 4354 590
rect 4253 525 4285 559
rect 4320 525 4354 559
rect 4253 494 4354 525
rect 310 415 400 425
rect 310 381 325 415
rect 359 381 400 415
rect 310 375 400 381
rect 1590 415 1680 425
rect 1590 381 1605 415
rect 1639 381 1680 415
rect 1590 375 1680 381
rect 2340 407 2410 425
rect 2340 373 2355 407
rect 2389 373 2410 407
rect 1066 339 1130 370
rect 2340 360 2410 373
rect 2865 415 2955 425
rect 2865 381 2885 415
rect 2919 381 2955 415
rect 2865 369 2955 381
rect 4150 415 4240 425
rect 4150 381 4165 415
rect 4199 381 4240 415
rect 4150 370 4240 381
rect 4900 407 4970 425
rect 4900 373 4915 407
rect 4949 373 4970 407
rect 4900 360 4970 373
rect 20 301 760 330
rect 20 300 634 301
rect 20 260 80 300
rect -80 247 80 260
rect -80 213 32 247
rect 66 213 80 247
rect -80 209 80 213
rect 160 247 220 260
rect 160 213 173 247
rect 207 213 220 247
rect 160 210 220 213
rect 20 200 80 209
rect 157 190 220 210
rect 579 247 640 260
rect 579 213 593 247
rect 627 213 640 247
rect 579 190 640 213
rect 690 247 760 301
rect 1066 305 1075 339
rect 1109 305 1130 339
rect 3620 339 3690 355
rect 1066 286 1130 305
rect 1300 300 2040 330
rect 690 213 710 247
rect 744 213 760 247
rect 690 200 760 213
rect 1300 247 1360 300
rect 1300 213 1312 247
rect 1346 213 1360 247
rect 1300 200 1360 213
rect 1440 247 1500 260
rect 1440 213 1453 247
rect 1487 213 1500 247
rect 1440 200 1500 213
rect 1860 247 1930 260
rect 1860 213 1873 247
rect 1907 213 1930 247
rect 157 160 640 190
rect 1440 170 1470 200
rect 1860 170 1930 213
rect 1980 247 2040 300
rect 1980 213 1990 247
rect 2024 213 2040 247
rect 1980 200 2040 213
rect 2580 300 3310 330
rect 2580 247 2640 300
rect 2580 213 2592 247
rect 2626 213 2640 247
rect 2580 200 2640 213
rect 2720 247 2780 260
rect 2720 213 2733 247
rect 2767 213 2780 247
rect 1440 141 1930 170
rect 1500 140 1930 141
rect 2720 170 2780 213
rect 3260 247 3310 300
rect 3620 305 3635 339
rect 3669 305 3690 339
rect 3620 290 3690 305
rect 3860 300 4600 330
rect 3260 213 3270 247
rect 3304 213 3310 247
rect 3260 200 3310 213
rect 3390 247 3450 260
rect 3390 213 3405 247
rect 3439 213 3450 247
rect 3390 170 3450 213
rect 3860 247 3920 300
rect 3860 213 3872 247
rect 3906 213 3920 247
rect 3860 199 3920 213
rect 4000 247 4060 260
rect 4430 259 4480 260
rect 4000 213 4013 247
rect 4047 213 4060 247
rect 2720 140 3450 170
rect 4000 170 4060 213
rect 4420 247 4480 259
rect 4420 213 4433 247
rect 4467 213 4480 247
rect 4420 170 4480 213
rect 4540 247 4600 300
rect 4540 213 4550 247
rect 4584 213 4600 247
rect 4540 200 4600 213
rect 4000 140 4480 170
rect 405 15 515 45
rect 405 -20 444 15
rect 480 -20 515 15
rect 405 -50 515 -20
rect 1144 15 1246 46
rect 1690 15 1796 46
rect 1144 -19 1174 15
rect 1210 -19 1246 15
rect 1686 -19 1725 15
rect 1760 -19 1796 15
rect 1144 -50 1246 -19
rect 1690 -50 1796 -19
rect 2424 15 2524 46
rect 2424 -19 2460 15
rect 2495 -19 2524 15
rect 2424 -50 2524 -19
rect 2973 15 3073 46
rect 2973 -19 3005 15
rect 3040 -19 3073 15
rect 2973 -50 3073 -19
rect 3706 15 3804 46
rect 3706 -19 3740 15
rect 3775 -19 3804 15
rect 3706 -50 3804 -19
rect 4252 15 4355 46
rect 4252 -19 4285 15
rect 4320 -19 4355 15
rect 4252 -50 4355 -19
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_0
timestamp 1691611044
transform 1 0 -42 0 1 -2
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_1
timestamp 1691611044
transform 1 0 1238 0 1 -2
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_2
timestamp 1691611044
transform 1 0 2518 0 1 -2
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  sky130_fd_sc_hd__and2_1_3
timestamp 1691611044
transform 1 0 3798 0 1 -2
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_0
timestamp 1691611044
transform 1 0 508 0 1 -2
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_1
timestamp 1691611044
transform 1 0 1788 0 1 -2
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_2
timestamp 1691611044
transform 1 0 3068 0 1 -2
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_3
timestamp 1691611044
transform 1 0 4348 0 1 -2
box -38 -48 682 592
<< labels >>
flabel metal1 0 260 0 260 1 FreeSans 320 0 0 0 A1
port 1 n
flabel metal1 1300 240 1300 240 1 FreeSans 320 0 0 0 A2
port 3 n
flabel viali 2610 240 2610 240 1 FreeSans 256 0 0 0 A3
port 5 n
flabel viali 3420 240 3420 240 1 FreeSans 192 0 0 0 B3
port 6 n
flabel viali 3888 240 3888 240 1 FreeSans 192 0 0 0 A4
port 7 n
flabel viali 610 240 610 240 1 FreeSans 192 0 0 0 B1
port 2 n
flabel viali 1890 242 1890 242 1 FreeSans 192 0 0 0 B2
port 4 n
flabel viali 4452 238 4452 238 1 FreeSans 192 0 0 0 B4
port 8 n
flabel viali 1090 330 1090 330 1 FreeSans 192 0 0 0 P1
port 10 n
flabel viali 340 405 340 405 1 FreeSans 128 0 0 0 G1
port 9 n
flabel viali 1620 405 1620 405 1 FreeSans 160 0 0 0 G2
port 11 n
flabel viali 2370 400 2370 400 1 FreeSans 128 0 0 0 P2
port 12 n
flabel viali 4930 400 4930 400 1 FreeSans 128 0 0 0 P4
port 16 n
flabel viali 3650 326 3650 326 1 FreeSans 256 0 0 0 P3
port 14 n
flabel viali 2900 400 2900 400 1 FreeSans 160 0 0 0 G3
port 13 n
flabel viali 4178 400 4178 400 1 FreeSans 160 0 0 0 G4
port 15 n
flabel viali s 96 0 96 0 1 FreeSans 160 0 0 0 GND
port 18 n
flabel viali 96 550 96 550 1 FreeSans 64 0 0 0 VDD
port 17 n
flabel nwell s 90 570 90 570 1 FreeSans 96 0 0 0 VPB
port 19 n
flabel pwell s 96 -34 96 -34 1 FreeSans 96 0 0 0 VNB
port 20 n
<< end >>
