magic
tech sky130A
magscale 1 2
timestamp 1703693701
<< nwell >>
rect -50 269 -47 590
rect 566 269 597 590
rect 1213 269 1238 590
rect 2726 269 2780 590
<< pwell >>
rect 523 56 634 211
rect 1173 56 1273 211
rect 1809 56 1902 203
rect 1982 56 2067 165
rect 2703 56 2810 211
<< locali >>
rect 537 535 564 569
rect 600 535 634 569
rect 1172 535 1210 569
rect 1245 535 1271 569
rect 1812 535 1840 569
rect 1875 535 1897 569
rect 1986 535 2010 569
rect 2045 535 2064 569
rect 2700 535 2736 569
rect 2771 535 2810 569
rect 1300 467 1335 470
rect 1300 435 1305 467
rect 1748 250 1782 257
rect 1748 223 1750 250
rect -10 135 50 150
rect -10 100 10 135
rect 44 100 50 135
rect 2630 145 2685 150
rect 2630 110 2640 145
rect 2675 110 2685 145
rect 2630 100 2685 110
rect -10 90 50 100
rect 527 -9 565 25
rect 600 -9 634 25
rect 1173 -9 1210 25
rect 1245 -9 1272 25
rect 1813 -9 1840 25
rect 1875 -9 1897 25
rect 1982 -9 2010 25
rect 2045 -9 2067 25
rect 2698 -9 2740 25
rect 2776 -9 2809 25
<< viali >>
rect 564 535 600 569
rect 1210 535 1245 569
rect 1840 535 1875 569
rect 2010 535 2045 569
rect 2736 535 2771 569
rect 1305 433 1339 467
rect 655 285 690 320
rect 212 223 246 257
rect 340 223 374 257
rect 468 223 502 257
rect 852 223 886 257
rect 980 223 1014 257
rect 1108 223 1142 257
rect 1492 223 1526 257
rect 1620 223 1654 257
rect 1750 215 1785 250
rect 2095 223 2129 257
rect 2241 223 2275 257
rect 2356 223 2392 258
rect 2456 223 2491 257
rect 2836 198 2871 233
rect 3027 223 3062 257
rect 3156 223 3190 257
rect 3284 223 3318 257
rect 10 100 44 135
rect 2640 110 2675 145
rect 565 -9 600 25
rect 1210 -9 1245 25
rect 1840 -9 1875 25
rect 2010 -9 2045 25
rect 2740 -9 2776 25
<< metal1 >>
rect 534 569 635 600
rect 534 535 564 569
rect 600 535 635 569
rect 534 504 635 535
rect 1175 569 1273 600
rect 1175 535 1210 569
rect 1245 535 1273 569
rect 1175 504 1273 535
rect 1818 569 1897 600
rect 1818 535 1840 569
rect 1875 535 1897 569
rect 1818 504 1897 535
rect 1987 569 2065 600
rect 1987 535 2010 569
rect 2045 535 2065 569
rect 1987 504 2065 535
rect 2698 569 2811 600
rect 2698 535 2736 569
rect 2771 535 2811 569
rect 2698 504 2811 535
rect 1285 467 3060 475
rect 1285 433 1305 467
rect 1339 445 3060 467
rect 1339 433 1345 445
rect 1285 420 1345 433
rect 470 360 2270 390
rect 470 280 500 360
rect 640 320 1660 330
rect 640 285 655 320
rect 690 300 1660 320
rect 690 285 710 300
rect 185 270 275 280
rect 185 200 195 270
rect 265 200 275 270
rect 185 190 275 200
rect 315 270 405 280
rect 315 200 325 270
rect 395 200 405 270
rect 315 190 405 200
rect 450 270 540 280
rect 640 275 710 285
rect 1610 270 1660 300
rect 2240 288 2270 360
rect 2216 278 2306 288
rect 3030 278 3060 445
rect 450 200 460 270
rect 530 200 540 270
rect 450 190 540 200
rect 830 260 910 270
rect 830 200 840 260
rect 900 200 910 260
rect 830 190 910 200
rect 970 257 1020 270
rect 970 223 980 257
rect 1014 223 1020 257
rect 970 150 1020 223
rect 1090 260 1170 270
rect 1090 200 1100 260
rect 1160 200 1170 260
rect 1090 190 1170 200
rect 1470 260 1550 270
rect 1470 205 1480 260
rect 1540 205 1550 260
rect 1610 257 1665 270
rect 1610 223 1620 257
rect 1654 223 1665 257
rect 1610 210 1665 223
rect 1725 260 1805 270
rect 1470 195 1550 205
rect 1725 205 1735 260
rect 1795 250 1805 260
rect 2081 257 2141 273
rect 2081 250 2095 257
rect 1795 223 2095 250
rect 2129 223 2141 257
rect 1795 220 2141 223
rect 1795 205 1805 220
rect 2081 208 2141 220
rect 2216 208 2226 278
rect 2296 208 2306 278
rect 2336 258 2406 268
rect 2336 223 2356 258
rect 2392 223 2406 258
rect 2336 210 2406 223
rect 2435 258 2520 270
rect 1725 195 1805 205
rect 2216 198 2306 208
rect -10 135 1020 150
rect -10 100 10 135
rect 44 120 1020 135
rect 1110 160 1140 190
rect 2355 160 2385 210
rect 2435 198 2446 258
rect 2506 198 2520 258
rect 3016 257 3076 278
rect 2435 185 2520 198
rect 2821 233 2885 248
rect 2821 198 2836 233
rect 2871 198 2885 233
rect 3016 223 3027 257
rect 3062 223 3076 257
rect 3016 205 3076 223
rect 3146 257 3196 273
rect 3146 223 3156 257
rect 3190 223 3196 257
rect 3146 210 3196 223
rect 3271 257 3336 273
rect 3271 223 3284 257
rect 3318 223 3336 257
rect 2821 173 2885 198
rect 1110 130 2385 160
rect 2625 145 2690 155
rect 3160 145 3190 210
rect 3271 208 3336 223
rect 44 100 59 120
rect 2625 110 2640 145
rect 2675 115 3190 145
rect 2675 110 2690 115
rect 2625 100 2690 110
rect -10 90 59 100
rect 533 25 634 56
rect 533 -9 565 25
rect 600 -9 634 25
rect 533 -40 634 -9
rect 1176 25 1272 56
rect 1176 -9 1210 25
rect 1245 -9 1272 25
rect 1176 -40 1272 -9
rect 1818 25 1899 56
rect 1818 -9 1840 25
rect 1875 -9 1899 25
rect 1818 -40 1899 -9
rect 1983 25 2068 56
rect 1983 -9 2010 25
rect 2045 -9 2068 25
rect 1983 -40 2068 -9
rect 2703 25 2810 56
rect 2703 -9 2740 25
rect 2776 -9 2810 25
rect 2703 -40 2810 -9
<< via1 >>
rect 195 257 265 270
rect 195 223 212 257
rect 212 223 246 257
rect 246 223 265 257
rect 195 200 265 223
rect 325 257 395 270
rect 325 223 340 257
rect 340 223 374 257
rect 374 223 395 257
rect 325 200 395 223
rect 460 257 530 270
rect 460 223 468 257
rect 468 223 502 257
rect 502 223 530 257
rect 460 200 530 223
rect 840 257 900 260
rect 840 223 852 257
rect 852 223 886 257
rect 886 223 900 257
rect 840 200 900 223
rect 1100 257 1160 260
rect 1100 223 1108 257
rect 1108 223 1142 257
rect 1142 223 1160 257
rect 1100 200 1160 223
rect 1480 257 1540 260
rect 1480 223 1492 257
rect 1492 223 1526 257
rect 1526 223 1540 257
rect 1480 205 1540 223
rect 1735 250 1795 260
rect 1735 215 1750 250
rect 1750 215 1785 250
rect 1785 215 1795 250
rect 1735 205 1795 215
rect 2226 257 2296 278
rect 2226 223 2241 257
rect 2241 223 2275 257
rect 2275 223 2296 257
rect 2226 208 2296 223
rect 2446 257 2506 258
rect 2446 223 2456 257
rect 2456 223 2491 257
rect 2491 223 2506 257
rect 2446 198 2506 223
<< metal2 >>
rect 185 270 275 280
rect 185 200 195 270
rect 265 200 275 270
rect 185 190 275 200
rect 315 270 405 280
rect 315 200 325 270
rect 395 200 405 270
rect 315 190 405 200
rect 450 270 540 280
rect 2216 278 2306 288
rect 450 200 460 270
rect 530 200 540 270
rect 450 190 540 200
rect 830 260 910 270
rect 830 200 840 260
rect 900 200 910 260
rect 830 190 910 200
rect 1090 260 1170 270
rect 1090 200 1100 260
rect 1160 200 1170 260
rect 1090 190 1170 200
rect 1470 260 1550 270
rect 1470 205 1480 260
rect 1540 205 1550 260
rect 1470 195 1550 205
rect 1725 260 1805 270
rect 1725 205 1735 260
rect 1795 205 1805 260
rect 1725 195 1805 205
rect 2216 208 2226 278
rect 2296 208 2306 278
rect 2216 198 2306 208
rect 2435 258 2520 270
rect 2435 198 2446 258
rect 2506 198 2520 258
rect 2435 185 2520 198
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_0
timestamp 1691611044
transform 1 0 -12 0 1 8
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_1
timestamp 1691611044
transform 1 0 628 0 1 8
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_2
timestamp 1691611044
transform 1 0 1268 0 1 8
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_3
timestamp 1691611044
transform 1 0 2804 0 1 8
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  sky130_fd_sc_hd__and4_1_0
timestamp 1691611044
transform 1 0 2064 0 1 8
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1691611044
transform 1 0 1896 0 1 8
box -38 -48 130 592
<< labels >>
flabel metal2 1130 270 1130 270 1 FreeSans 128 0 0 0 P3
port 6 n
flabel metal1 870 270 870 270 1 FreeSans 128 0 0 0 G3
port 7 n
flabel metal1 1510 270 1510 270 1 FreeSans 128 0 0 0 G4
port 9 n
flabel metal2 490 270 490 270 1 FreeSans 128 0 0 0 P2
port 4 n
flabel metal1 350 270 350 270 1 FreeSans 128 0 0 0 G1
port 3 n
flabel viali 230 225 230 225 1 FreeSans 128 0 0 0 G2
port 5 n
flabel metal1 3306 268 3306 268 1 FreeSans 128 0 0 0 CI
port 1 n
flabel metal1 2826 213 2826 213 1 FreeSans 128 0 0 0 CO
port 10 n
flabel via1 1765 245 1765 245 1 FreeSans 320 0 0 0 P4
port 8 n
flabel via1 2465 250 2465 250 1 FreeSans 160 0 0 0 P1
port 2 n
flabel space 10 575 10 575 1 FreeSans 320 0 0 0 VDD
port 11 n
flabel space 0 5 0 5 1 FreeSans 320 0 0 0 GND
port 12 n
flabel locali s 1935 345 1935 345 1 FreeSans 320 0 0 0 VPB
port 13 n
flabel locali s 1940 130 1940 130 1 FreeSans 320 0 0 0 VNB
port 14 n
<< end >>
