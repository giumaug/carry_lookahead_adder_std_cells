magic
tech sky130A
magscale 1 2
timestamp 1703239092
<< locali >>
rect -140 599 -130 633
rect -95 599 -41 633
rect -5 599 21 633
rect 5202 55 5240 89
rect 5275 55 5330 89
rect 5365 55 5420 89
rect 5455 55 5510 89
rect 5545 55 5610 89
rect 5645 55 5685 89
rect -140 -742 -130 -708
rect -95 -742 -45 -708
rect -10 -742 22 -708
rect 3383 -1286 3415 -1252
rect 3450 -1286 3505 -1252
rect 3540 -1286 3595 -1252
rect 3630 -1286 3685 -1252
rect 3720 -1286 3775 -1252
rect 3810 -1286 3865 -1252
rect 3900 -1286 3955 -1252
rect 3990 -1286 4045 -1252
rect 4080 -1286 4135 -1252
rect 4170 -1286 4225 -1252
rect 4260 -1286 4315 -1252
rect 4350 -1286 4405 -1252
rect 4440 -1286 4495 -1252
rect 4530 -1286 4585 -1252
rect 4620 -1286 4675 -1252
rect 4710 -1286 4765 -1252
rect 4800 -1286 4855 -1252
rect 4890 -1286 4945 -1252
rect 4980 -1286 5035 -1252
rect 5070 -1286 5125 -1252
rect 5160 -1286 5215 -1252
rect 5250 -1286 5305 -1252
rect 5340 -1286 5395 -1252
rect 5430 -1286 5485 -1252
rect 5520 -1286 5575 -1252
rect 5610 -1286 5660 -1252
rect -140 -1525 -130 -1491
rect -95 -1525 -45 -1491
rect -10 -1525 22 -1491
rect 5547 -2069 5575 -2035
rect 5610 -2069 5660 -2035
<< viali >>
rect -130 599 -95 633
rect -41 599 -5 633
rect 5240 55 5275 89
rect 5330 55 5365 89
rect 5420 55 5455 89
rect 5510 55 5545 89
rect 5610 55 5645 89
rect -130 -742 -95 -708
rect -45 -742 -10 -708
rect 3415 -1286 3450 -1252
rect 3505 -1286 3540 -1252
rect 3595 -1286 3630 -1252
rect 3685 -1286 3720 -1252
rect 3775 -1286 3810 -1252
rect 3865 -1286 3900 -1252
rect 3955 -1286 3990 -1252
rect 4045 -1286 4080 -1252
rect 4135 -1286 4170 -1252
rect 4225 -1286 4260 -1252
rect 4315 -1286 4350 -1252
rect 4405 -1286 4440 -1252
rect 4495 -1286 4530 -1252
rect 4585 -1286 4620 -1252
rect 4675 -1286 4710 -1252
rect 4765 -1286 4800 -1252
rect 4855 -1286 4890 -1252
rect 4945 -1286 4980 -1252
rect 5035 -1286 5070 -1252
rect 5125 -1286 5160 -1252
rect 5215 -1286 5250 -1252
rect 5305 -1286 5340 -1252
rect 5395 -1286 5430 -1252
rect 5485 -1286 5520 -1252
rect 5575 -1286 5610 -1252
rect 5660 -1286 5695 -1252
rect -130 -1525 -95 -1491
rect -45 -1525 -10 -1491
rect 5575 -2069 5610 -2035
rect 5660 -2069 5695 -2035
<< metal1 >>
rect 3290 1445 3370 1455
rect 3290 1430 3300 1445
rect -140 1400 3300 1430
rect 3290 1385 3300 1400
rect 3360 1385 3370 1445
rect 3290 1375 3370 1385
rect 4630 1360 4710 1370
rect 4630 1345 4640 1360
rect -140 1315 4640 1345
rect 4630 1300 4640 1315
rect 4700 1300 4710 1360
rect 4630 1290 4710 1300
rect 4065 1275 4145 1285
rect 4065 1260 4075 1275
rect -140 1230 4075 1260
rect 4065 1215 4075 1230
rect 4135 1215 4145 1275
rect 4065 1205 4145 1215
rect 3600 1190 3680 1200
rect 3600 1175 3610 1190
rect -140 1145 3610 1175
rect 3600 1130 3610 1145
rect 3670 1130 3680 1190
rect 3600 1120 3680 1130
rect 2785 1105 2865 1115
rect 2785 1090 2795 1105
rect -140 1060 2795 1090
rect 2785 1045 2795 1060
rect 2855 1045 2865 1105
rect 2785 1035 2865 1045
rect 1910 1020 1990 1030
rect 1910 1005 1920 1020
rect -140 975 1920 1005
rect 1910 960 1920 975
rect 1980 960 1990 1020
rect 1910 950 1990 960
rect 1350 935 1425 945
rect 1350 920 1360 935
rect -140 890 1360 920
rect 1350 875 1360 890
rect 1415 875 1425 935
rect 1350 865 1425 875
rect 635 850 715 860
rect 635 835 645 850
rect -140 805 645 835
rect 635 790 645 805
rect 705 790 715 850
rect 635 780 715 790
rect 70 765 150 775
rect 70 750 80 765
rect -140 720 80 750
rect 70 705 80 720
rect 140 705 150 765
rect 70 695 150 705
rect -140 650 23 664
rect -140 633 -100 650
rect -40 633 23 650
rect -140 599 -130 633
rect -5 599 23 633
rect -140 590 -100 599
rect -40 590 23 599
rect -140 568 23 590
rect 360 510 440 520
rect 360 450 370 510
rect 430 450 440 510
rect 360 440 440 450
rect 1640 515 1720 525
rect 1640 455 1650 515
rect 1710 455 1720 515
rect 1640 445 1720 455
rect 2390 500 2470 510
rect 1110 435 1190 445
rect 1110 375 1120 435
rect 1180 375 1190 435
rect 2390 440 2400 500
rect 2460 440 2470 500
rect 2390 430 2470 440
rect 3080 505 3160 515
rect 3080 445 3090 505
rect 3150 445 3160 505
rect 3080 435 3160 445
rect 4360 510 4435 520
rect 4360 450 4370 510
rect 4425 450 4435 510
rect 4360 440 4435 450
rect 5110 495 5190 505
rect 3830 430 3910 440
rect 1110 365 1190 375
rect 3830 370 3840 430
rect 3900 370 3910 430
rect 5110 435 5120 495
rect 5180 435 5190 495
rect 5110 425 5190 435
rect 3830 360 3910 370
rect 70 335 150 345
rect 70 275 80 335
rect 140 275 150 335
rect 70 265 150 275
rect 635 335 715 345
rect 635 275 645 335
rect 705 275 715 335
rect 635 260 715 275
rect 1350 335 1430 345
rect 1350 275 1360 335
rect 1420 275 1430 335
rect 1350 265 1430 275
rect 1910 335 1990 345
rect 1910 275 1920 335
rect 1980 275 1990 335
rect 1910 265 1990 275
rect 2785 330 2865 340
rect 2785 270 2795 330
rect 2855 270 2865 330
rect 1910 230 1920 265
rect 2785 260 2865 270
rect 3600 330 3680 340
rect 3600 270 3610 330
rect 3670 270 3680 330
rect 3600 260 3680 270
rect 4065 330 4145 340
rect 4065 270 4075 330
rect 4135 270 4145 330
rect 4065 260 4145 270
rect 4630 330 4710 340
rect 4630 270 4640 330
rect 4700 270 4710 330
rect 4630 260 4710 270
rect 3600 225 3615 260
rect 4630 225 4645 260
rect 5205 100 5705 120
rect 5205 89 5605 100
rect 5205 55 5240 89
rect 5275 55 5330 89
rect 5365 55 5420 89
rect 5455 55 5510 89
rect 5545 55 5605 89
rect 5205 40 5605 55
rect 5665 40 5705 100
rect 5205 25 5705 40
rect 95 -15 175 -5
rect 95 -30 105 -15
rect 50 -60 105 -30
rect 95 -75 105 -60
rect 165 -30 175 -15
rect 360 -15 440 -5
rect 360 -30 370 -15
rect 165 -60 370 -30
rect 165 -75 175 -60
rect 95 -85 175 -75
rect 360 -75 370 -60
rect 430 -75 440 -15
rect 360 -85 440 -75
rect 860 -15 940 -5
rect 860 -75 870 -15
rect 930 -30 940 -15
rect 1375 -15 1455 -5
rect 1375 -30 1385 -15
rect 930 -60 1385 -30
rect 930 -75 940 -60
rect 860 -85 940 -75
rect 1375 -75 1385 -60
rect 1445 -30 1455 -15
rect 3080 -15 3160 -5
rect 3080 -30 3090 -15
rect 1445 -60 3090 -30
rect 1445 -75 1455 -60
rect 1375 -85 1455 -75
rect 3080 -75 3090 -60
rect 3150 -75 3160 -15
rect 3080 -85 3160 -75
rect 220 -100 300 -90
rect 220 -115 230 -100
rect 120 -145 230 -115
rect 220 -160 230 -145
rect 290 -115 300 -100
rect 750 -100 830 -90
rect 750 -115 760 -100
rect 290 -145 760 -115
rect 290 -160 300 -145
rect 220 -170 300 -160
rect 750 -160 760 -145
rect 820 -115 830 -100
rect 1640 -100 1720 -90
rect 1640 -115 1650 -100
rect 820 -145 1650 -115
rect 820 -160 830 -145
rect 750 -170 830 -160
rect 1640 -160 1650 -145
rect 1710 -160 1720 -100
rect 1640 -170 1720 -160
rect 475 -185 555 -175
rect 475 -245 485 -185
rect 545 -200 555 -185
rect 1220 -185 1300 -175
rect 1220 -200 1230 -185
rect 545 -230 1230 -200
rect 545 -245 555 -230
rect 475 -255 555 -245
rect 1220 -245 1230 -230
rect 1290 -200 1300 -185
rect 2390 -185 2470 -175
rect 2390 -200 2400 -185
rect 1290 -230 2400 -200
rect 1290 -245 1300 -230
rect 1220 -255 1300 -245
rect 2390 -245 2400 -230
rect 2460 -245 2470 -185
rect 2390 -255 2470 -245
rect 575 -295 655 -285
rect 575 -355 585 -295
rect 645 -310 655 -295
rect 1110 -295 1190 -285
rect 1110 -310 1120 -295
rect 645 -340 1120 -310
rect 645 -355 655 -340
rect 575 -365 655 -355
rect 1110 -355 1120 -340
rect 1180 -310 1190 -295
rect 2470 -295 2550 -285
rect 2470 -310 2480 -295
rect 1180 -340 2480 -310
rect 1180 -355 1190 -340
rect 1110 -365 1190 -355
rect 2470 -355 2480 -340
rect 2540 -355 2550 -295
rect 2470 -365 2550 -355
rect 1115 -405 1195 -395
rect 1115 -465 1125 -405
rect 1185 -420 1195 -405
rect 1900 -405 1980 -395
rect 1900 -420 1910 -405
rect 1185 -450 1910 -420
rect 1185 -465 1195 -450
rect 1115 -475 1195 -465
rect 1900 -465 1910 -450
rect 1970 -420 1980 -405
rect 3830 -405 3910 -395
rect 3830 -420 3840 -405
rect 1970 -450 3840 -420
rect 1970 -465 1980 -450
rect 1900 -475 1980 -465
rect 3830 -465 3840 -450
rect 3900 -465 3910 -405
rect 3830 -475 3910 -465
rect 1500 -490 1580 -480
rect 1500 -550 1510 -490
rect 1570 -505 1580 -490
rect 2125 -490 2205 -480
rect 2125 -505 2135 -490
rect 1570 -535 2135 -505
rect 1570 -550 1580 -535
rect 1500 -560 1580 -550
rect 2125 -550 2135 -535
rect 2195 -505 2205 -490
rect 2380 -490 2460 -480
rect 2380 -505 2390 -490
rect 2195 -535 2390 -505
rect 2195 -550 2205 -535
rect 2125 -560 2205 -550
rect 2380 -550 2390 -535
rect 2450 -505 2460 -490
rect 4360 -490 4440 -480
rect 4360 -505 4370 -490
rect 2450 -535 4370 -505
rect 2450 -550 2460 -535
rect 2380 -560 2460 -550
rect 4360 -550 4370 -535
rect 4430 -550 4440 -490
rect 4360 -560 4440 -550
rect 1760 -575 1840 -565
rect 1760 -630 1770 -575
rect 1830 -590 1840 -575
rect 5110 -575 5190 -565
rect 5110 -590 5120 -575
rect 1830 -620 5120 -590
rect 1830 -630 1840 -620
rect 1760 -640 1840 -630
rect 5110 -635 5120 -620
rect 5180 -635 5190 -575
rect 5110 -645 5190 -635
rect -140 -695 22 -678
rect -140 -708 -100 -695
rect -40 -708 22 -695
rect -140 -742 -130 -708
rect -10 -742 22 -708
rect -140 -755 -100 -742
rect -40 -755 22 -742
rect -140 -773 22 -755
rect 3295 -1005 3375 -995
rect 1115 -1080 1195 -1005
rect 3295 -1065 3305 -1005
rect 3365 -1065 3375 -1005
rect 3295 -1075 3375 -1065
rect 1115 -1085 1120 -1080
rect 1140 -1085 1195 -1080
rect 3380 -1240 5705 -1221
rect 3380 -1252 5605 -1240
rect 5665 -1252 5705 -1240
rect 3380 -1286 3415 -1252
rect 3450 -1286 3505 -1252
rect 3540 -1286 3595 -1252
rect 3630 -1286 3685 -1252
rect 3720 -1286 3775 -1252
rect 3810 -1286 3865 -1252
rect 3900 -1286 3955 -1252
rect 3990 -1286 4045 -1252
rect 4080 -1286 4135 -1252
rect 4170 -1286 4225 -1252
rect 4260 -1286 4315 -1252
rect 4350 -1286 4405 -1252
rect 4440 -1286 4495 -1252
rect 4530 -1286 4585 -1252
rect 4620 -1286 4675 -1252
rect 4710 -1286 4765 -1252
rect 4800 -1286 4855 -1252
rect 4890 -1286 4945 -1252
rect 4980 -1286 5035 -1252
rect 5070 -1286 5125 -1252
rect 5160 -1286 5215 -1252
rect 5250 -1286 5305 -1252
rect 5340 -1286 5395 -1252
rect 5430 -1286 5485 -1252
rect 5520 -1286 5575 -1252
rect 5695 -1286 5705 -1252
rect 3380 -1300 5605 -1286
rect 5665 -1300 5705 -1286
rect 3380 -1317 5705 -1300
rect 345 -1360 425 -1350
rect 345 -1420 355 -1360
rect 415 -1375 425 -1360
rect 3295 -1360 3375 -1350
rect 3295 -1375 3305 -1360
rect 415 -1405 3305 -1375
rect 415 -1420 425 -1405
rect 345 -1430 425 -1420
rect 3295 -1420 3305 -1405
rect 3365 -1420 3375 -1360
rect 3295 -1430 3375 -1420
rect -140 -1475 29 -1460
rect -140 -1491 -100 -1475
rect -40 -1491 29 -1475
rect -140 -1525 -130 -1491
rect -10 -1525 29 -1491
rect -140 -1535 -100 -1525
rect -40 -1535 29 -1525
rect -140 -1556 29 -1535
rect 1745 -1599 1825 -1589
rect 1745 -1659 1755 -1599
rect 1815 -1614 1825 -1599
rect 1900 -1599 1980 -1589
rect 1900 -1614 1910 -1599
rect 1815 -1644 1910 -1614
rect 1815 -1659 1825 -1644
rect 1745 -1669 1825 -1659
rect 1900 -1659 1910 -1644
rect 1970 -1659 1980 -1599
rect 1900 -1669 1980 -1659
rect 5544 -2025 5705 -2004
rect 5544 -2035 5605 -2025
rect 5665 -2035 5705 -2025
rect 5544 -2069 5575 -2035
rect 5695 -2069 5705 -2035
rect 5544 -2085 5605 -2069
rect 5665 -2085 5705 -2069
rect 5544 -2100 5705 -2085
rect 3265 -2155 3345 -2130
rect 3265 -2185 5705 -2155
rect 3265 -2210 3345 -2185
rect 3990 -2225 4070 -2215
rect 3990 -2285 4000 -2225
rect 4060 -2240 4070 -2225
rect 4060 -2270 5705 -2240
rect 4060 -2285 4070 -2270
rect 3990 -2295 4070 -2285
rect 4720 -2310 4800 -2300
rect 4720 -2370 4730 -2310
rect 4790 -2325 4800 -2310
rect 4790 -2355 5705 -2325
rect 4790 -2370 4800 -2355
rect 4720 -2380 4800 -2370
rect 5450 -2395 5530 -2385
rect 5450 -2455 5460 -2395
rect 5520 -2410 5530 -2395
rect 5520 -2440 5705 -2410
rect 5520 -2455 5530 -2440
rect 5450 -2465 5530 -2455
rect 1930 -2650 2010 -2640
rect 1930 -2710 1940 -2650
rect 2000 -2665 2010 -2650
rect 2000 -2695 5705 -2665
rect 2000 -2710 2010 -2695
rect 1930 -2720 2010 -2710
<< via1 >>
rect 3300 1385 3360 1445
rect 4640 1300 4700 1360
rect 4075 1215 4135 1275
rect 3610 1130 3670 1190
rect 2795 1045 2855 1105
rect 1920 960 1980 1020
rect 1360 875 1415 935
rect 645 790 705 850
rect 80 705 140 765
rect -100 633 -40 650
rect -100 599 -95 633
rect -95 599 -41 633
rect -41 599 -40 633
rect -100 590 -40 599
rect 370 450 430 510
rect 1650 455 1710 515
rect 1120 375 1180 435
rect 2400 440 2460 500
rect 3090 445 3150 505
rect 4370 450 4425 510
rect 3840 370 3900 430
rect 5120 435 5180 495
rect 80 275 140 335
rect 645 275 705 335
rect 1360 275 1420 335
rect 1920 275 1980 335
rect 2795 270 2855 330
rect 3610 270 3670 330
rect 4075 270 4135 330
rect 4640 270 4700 330
rect 5605 89 5665 100
rect 5605 55 5610 89
rect 5610 55 5645 89
rect 5645 55 5665 89
rect 5605 40 5665 55
rect 105 -75 165 -15
rect 370 -75 430 -15
rect 870 -75 930 -15
rect 1385 -75 1445 -15
rect 3090 -75 3150 -15
rect 230 -160 290 -100
rect 760 -160 820 -100
rect 1650 -160 1710 -100
rect 485 -245 545 -185
rect 1230 -245 1290 -185
rect 2400 -245 2460 -185
rect 585 -355 645 -295
rect 1120 -355 1180 -295
rect 2480 -355 2540 -295
rect 1125 -465 1185 -405
rect 1910 -465 1970 -405
rect 3840 -465 3900 -405
rect 1510 -550 1570 -490
rect 2135 -550 2195 -490
rect 2390 -550 2450 -490
rect 4370 -550 4430 -490
rect 1770 -630 1830 -575
rect 5120 -635 5180 -575
rect -100 -708 -40 -695
rect -100 -742 -95 -708
rect -95 -742 -45 -708
rect -45 -742 -40 -708
rect -100 -755 -40 -742
rect 3305 -1065 3365 -1005
rect 5605 -1252 5665 -1240
rect 5605 -1286 5610 -1252
rect 5610 -1286 5660 -1252
rect 5660 -1286 5665 -1252
rect 5605 -1300 5665 -1286
rect 355 -1420 415 -1360
rect 3305 -1420 3365 -1360
rect -100 -1491 -40 -1475
rect -100 -1525 -95 -1491
rect -95 -1525 -45 -1491
rect -45 -1525 -40 -1491
rect -100 -1535 -40 -1525
rect 1755 -1659 1815 -1599
rect 1910 -1659 1970 -1599
rect 5605 -2035 5665 -2025
rect 5605 -2069 5610 -2035
rect 5610 -2069 5660 -2035
rect 5660 -2069 5665 -2035
rect 5605 -2085 5665 -2069
rect 4000 -2285 4060 -2225
rect 4730 -2370 4790 -2310
rect 5460 -2455 5520 -2395
rect 1940 -2710 2000 -2650
<< metal2 >>
rect 3290 1445 3370 1455
rect 3290 1385 3300 1445
rect 3360 1385 3370 1445
rect 3290 1375 3370 1385
rect 2785 1105 2865 1115
rect 2785 1045 2795 1105
rect 2855 1045 2865 1105
rect 2785 1035 2865 1045
rect 1910 1020 1990 1030
rect 1910 960 1920 1020
rect 1980 960 1990 1020
rect 1910 950 1990 960
rect 1350 935 1425 945
rect 1350 875 1360 935
rect 1415 875 1425 935
rect 1350 865 1425 875
rect 635 850 715 860
rect 635 790 645 850
rect 705 790 715 850
rect 635 780 715 790
rect 70 765 150 775
rect 70 705 80 765
rect 140 705 150 765
rect 70 695 150 705
rect -120 650 -20 670
rect -120 590 -100 650
rect -40 590 -20 650
rect -120 -695 -20 590
rect 95 345 125 695
rect 360 510 440 520
rect 360 450 370 510
rect 430 450 440 510
rect 360 440 440 450
rect 70 335 150 345
rect 70 275 80 335
rect 140 275 150 335
rect 70 265 150 275
rect 385 -5 415 440
rect 660 345 690 780
rect 1110 435 1190 445
rect 1110 375 1120 435
rect 1180 375 1190 435
rect 1110 365 1190 375
rect 635 335 715 345
rect 635 275 645 335
rect 705 275 715 335
rect 635 265 715 275
rect 95 -15 175 -5
rect 95 -75 105 -15
rect 165 -75 175 -15
rect 95 -85 175 -75
rect 360 -15 440 -5
rect 360 -75 370 -15
rect 430 -75 440 -15
rect 360 -85 440 -75
rect 860 -15 940 -5
rect 860 -75 870 -15
rect 930 -75 940 -15
rect 860 -85 940 -75
rect -120 -755 -100 -695
rect -40 -755 -20 -695
rect -120 -1475 -20 -755
rect -120 -1535 -100 -1475
rect -40 -1535 -20 -1475
rect -120 -1556 -20 -1535
rect 120 -1804 150 -85
rect 220 -100 300 -90
rect 220 -160 230 -100
rect 290 -160 300 -100
rect 220 -170 300 -160
rect 245 -1010 275 -170
rect 370 -1010 400 -85
rect 750 -100 830 -90
rect 750 -160 760 -100
rect 820 -160 830 -100
rect 750 -170 830 -160
rect 475 -185 555 -175
rect 475 -245 485 -185
rect 545 -245 555 -185
rect 475 -255 555 -245
rect 500 -1010 530 -255
rect 575 -295 655 -285
rect 575 -355 585 -295
rect 645 -355 655 -295
rect 575 -365 655 -355
rect 215 -1050 225 -1020
rect 550 -1050 560 -1020
rect 245 -1085 275 -1075
rect 370 -1085 400 -1075
rect 500 -1085 530 -1070
rect 345 -1360 425 -1350
rect 345 -1420 355 -1360
rect 415 -1420 425 -1360
rect 345 -1430 425 -1420
rect 370 -1800 400 -1430
rect 600 -1799 630 -365
rect 120 -1834 225 -1804
rect 560 -1829 630 -1799
rect 775 -1804 805 -170
rect 885 -1015 915 -85
rect 1135 -285 1165 365
rect 1375 345 1405 865
rect 1640 515 1720 525
rect 1640 455 1650 515
rect 1710 455 1720 515
rect 1640 445 1720 455
rect 1350 335 1430 345
rect 1350 275 1360 335
rect 1420 275 1430 335
rect 1350 265 1430 275
rect 1375 -15 1455 -5
rect 1375 -75 1385 -15
rect 1445 -75 1455 -15
rect 1375 -85 1455 -75
rect 1220 -185 1300 -175
rect 1220 -245 1230 -185
rect 1290 -245 1300 -185
rect 1220 -255 1300 -245
rect 1110 -295 1190 -285
rect 1110 -355 1120 -295
rect 1180 -355 1190 -295
rect 1110 -365 1190 -355
rect 1115 -405 1195 -395
rect 1115 -465 1125 -405
rect 1185 -465 1195 -405
rect 1115 -475 1195 -465
rect 1140 -1005 1170 -475
rect 885 -1085 915 -1060
rect 1115 -1085 1195 -1005
rect 1140 -1090 1170 -1085
rect 1245 -1804 1275 -255
rect 775 -1834 860 -1804
rect 1190 -1834 1275 -1804
rect 1400 -1804 1430 -85
rect 1665 -90 1695 445
rect 1935 345 1965 950
rect 2390 500 2470 510
rect 2390 440 2400 500
rect 2460 440 2470 500
rect 2390 430 2470 440
rect 1910 335 1990 345
rect 1910 275 1920 335
rect 1980 275 1990 335
rect 1910 265 1990 275
rect 1640 -100 1720 -90
rect 1640 -160 1650 -100
rect 1710 -160 1720 -100
rect 1640 -170 1720 -160
rect 2415 -175 2445 430
rect 2810 340 2840 1035
rect 3080 505 3160 515
rect 3080 445 3090 505
rect 3150 445 3160 505
rect 3080 435 3160 445
rect 2785 330 2865 340
rect 2785 270 2795 330
rect 2855 270 2865 330
rect 2785 260 2865 270
rect 3105 -5 3135 435
rect 3080 -15 3160 -5
rect 3080 -75 3090 -15
rect 3150 -75 3160 -15
rect 3080 -85 3160 -75
rect 2390 -185 2470 -175
rect 2390 -245 2400 -185
rect 2460 -245 2470 -185
rect 2390 -255 2470 -245
rect 2470 -295 2550 -285
rect 2470 -355 2480 -295
rect 2540 -355 2550 -295
rect 2470 -365 2550 -355
rect 1900 -405 1980 -395
rect 1900 -465 1910 -405
rect 1970 -465 1980 -405
rect 1900 -475 1980 -465
rect 1500 -490 1580 -480
rect 1500 -550 1510 -490
rect 1570 -550 1580 -490
rect 1500 -560 1580 -550
rect 1525 -1015 1555 -560
rect 1760 -575 1840 -565
rect 1760 -630 1770 -575
rect 1830 -630 1840 -575
rect 1760 -640 1840 -630
rect 1785 -1015 1815 -640
rect 1525 -1080 1555 -1060
rect 1785 -1080 1815 -1065
rect 1925 -1589 1955 -475
rect 2125 -490 2205 -480
rect 2125 -550 2135 -490
rect 2195 -550 2205 -490
rect 2125 -560 2205 -550
rect 2380 -490 2460 -480
rect 2380 -550 2390 -490
rect 2450 -550 2460 -490
rect 2380 -560 2460 -550
rect 1745 -1599 1825 -1589
rect 1745 -1659 1755 -1599
rect 1815 -1659 1825 -1599
rect 1745 -1669 1825 -1659
rect 1900 -1599 1980 -1589
rect 1900 -1659 1910 -1599
rect 1970 -1659 1980 -1599
rect 1900 -1669 1980 -1659
rect 1770 -1799 1800 -1669
rect 2150 -1794 2180 -560
rect 2405 -1799 2435 -560
rect 2490 -1045 2520 -365
rect 3315 -995 3345 1375
rect 4630 1360 4710 1370
rect 4630 1300 4640 1360
rect 4700 1300 4710 1360
rect 4630 1290 4710 1300
rect 4065 1275 4145 1285
rect 4065 1215 4075 1275
rect 4135 1215 4145 1275
rect 4065 1205 4145 1215
rect 3600 1190 3680 1200
rect 3600 1130 3610 1190
rect 3670 1130 3680 1190
rect 3600 1120 3680 1130
rect 3625 340 3655 1120
rect 3830 430 3910 440
rect 3830 370 3840 430
rect 3900 370 3910 430
rect 3830 360 3910 370
rect 3600 330 3680 340
rect 3600 270 3610 330
rect 3670 270 3680 330
rect 3600 260 3680 270
rect 3855 -395 3885 360
rect 4090 340 4120 1205
rect 4360 510 4435 520
rect 4360 450 4370 510
rect 4425 450 4435 510
rect 4360 440 4435 450
rect 4065 330 4145 340
rect 4065 270 4075 330
rect 4135 270 4145 330
rect 4065 260 4145 270
rect 3830 -405 3910 -395
rect 3830 -465 3840 -405
rect 3900 -465 3910 -405
rect 3830 -475 3910 -465
rect 4385 -480 4415 440
rect 4655 340 4685 1290
rect 5110 495 5190 505
rect 5110 435 5120 495
rect 5180 435 5190 495
rect 5110 425 5190 435
rect 4630 330 4710 340
rect 4630 270 4640 330
rect 4700 270 4710 330
rect 4630 260 4710 270
rect 4360 -490 4440 -480
rect 4360 -550 4370 -490
rect 4430 -550 4440 -490
rect 4360 -560 4440 -550
rect 5135 -565 5165 425
rect 5585 100 5685 120
rect 5585 40 5605 100
rect 5665 40 5685 100
rect 5110 -575 5190 -565
rect 5110 -635 5120 -575
rect 5180 -635 5190 -575
rect 5110 -645 5190 -635
rect 3295 -1005 3375 -995
rect 2490 -1090 2520 -1060
rect 3295 -1065 3305 -1005
rect 3365 -1065 3375 -1005
rect 3295 -1075 3375 -1065
rect 3320 -1350 3350 -1075
rect 5585 -1240 5685 40
rect 5585 -1300 5605 -1240
rect 5665 -1300 5685 -1240
rect 3295 -1360 3375 -1350
rect 3295 -1420 3305 -1360
rect 3365 -1420 3375 -1360
rect 3295 -1430 3375 -1420
rect 1400 -1834 1495 -1804
rect 1955 -2640 1985 -1830
rect 3290 -2130 3320 -1760
rect 3265 -2210 3345 -2130
rect 4015 -2215 4045 -1745
rect 3990 -2225 4070 -2215
rect 3990 -2285 4000 -2225
rect 4060 -2285 4070 -2225
rect 3990 -2295 4070 -2285
rect 4745 -2300 4775 -1755
rect 4720 -2310 4800 -2300
rect 4720 -2370 4730 -2310
rect 4790 -2370 4800 -2310
rect 4720 -2380 4800 -2370
rect 5475 -2385 5505 -1745
rect 5585 -2025 5685 -1300
rect 5585 -2085 5605 -2025
rect 5665 -2085 5685 -2025
rect 5585 -2100 5685 -2085
rect 5450 -2395 5530 -2385
rect 5450 -2455 5460 -2395
rect 5520 -2455 5530 -2395
rect 5450 -2465 5530 -2455
rect 1930 -2650 2010 -2640
rect 1930 -2710 1940 -2650
rect 2000 -2710 2010 -2650
rect 1930 -2720 2010 -2710
use adder_1  adder_1_0
timestamp 1700079872
transform 1 0 60 0 1 74
box -80 -50 5188 590
use adder_2  adder_2_0
timestamp 1700046346
transform 1 0 30 0 1 -1277
box -50 -40 3394 600
use adder_3  adder_3_0
timestamp 1699994886
transform 1 0 25 0 1 -2055
box -45 -580 5561 595
<< labels >>
flabel metal1 20 735 20 735 1 FreeSans 160 0 0 0 A1
port 1 n
flabel metal1 25 820 25 820 1 FreeSans 160 0 0 0 B1
port 2 n
flabel metal1 25 905 25 905 1 FreeSans 160 0 0 0 A2
port 3 n
flabel metal1 25 990 25 990 1 FreeSans 160 0 0 0 B2
port 4 n
flabel metal1 25 1075 25 1075 1 FreeSans 160 0 0 0 A3
port 5 n
flabel metal1 25 1160 25 1160 1 FreeSans 160 0 0 0 B3
port 6 n
flabel metal1 25 1245 25 1245 1 FreeSans 160 0 0 0 A4
port 7 n
flabel metal1 25 1330 25 1330 1 FreeSans 160 0 0 0 B4
port 8 n
flabel metal1 25 1415 25 1415 1 FreeSans 160 0 0 0 CI
port 9 n
flabel metal1 5700 -2170 5700 -2170 7 FreeSans 160 0 0 0 S1
port 10 w
flabel metal1 5700 -2255 5700 -2255 7 FreeSans 160 0 0 0 S2
port 11 w
flabel metal1 5700 -2340 5700 -2340 7 FreeSans 160 0 0 0 S3
port 12 w
flabel metal1 5700 -2425 5700 -2425 7 FreeSans 160 0 0 0 S4
port 13 w
flabel metal1 5700 -2680 5700 -2680 7 FreeSans 160 0 0 0 CO
port 14 w
flabel via1 -75 619 -75 619 1 FreeSans 128 0 0 0 VDD
port 15 n
flabel via1 5635 -2055 5635 -2055 1 FreeSans 128 0 0 0 GND
port 16 n
<< end >>
