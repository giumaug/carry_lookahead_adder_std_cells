magic
tech sky130A
magscale 1 2
timestamp 1699994886
<< nwell >>
rect 570 264 596 585
rect 1212 264 1231 585
rect 1851 264 1862 585
rect 3366 264 3388 585
rect 4091 264 4114 585
rect 4824 264 4850 585
<< pwell >>
rect 537 51 634 206
rect 1170 51 1269 206
rect 1808 51 1903 206
rect 2436 51 2534 198
rect 2601 51 2708 198
rect 3331 51 3434 205
rect 4053 51 4162 206
rect 4782 51 4892 206
<< locali >>
rect 542 530 575 564
rect 610 530 636 564
rect 1171 530 1205 564
rect 1240 530 1269 564
rect 1810 530 1840 564
rect 1875 530 1903 564
rect 2437 530 2470 564
rect 2505 530 2529 564
rect 2603 530 2640 564
rect 2675 530 2699 564
rect 3334 530 3361 564
rect 3396 530 3428 564
rect 4053 530 4091 564
rect 4126 530 4155 564
rect 4783 530 4816 564
rect 4851 530 4885 564
rect 665 460 699 462
rect 660 430 699 460
rect 690 428 699 430
rect 1300 428 1334 462
rect 690 425 695 428
rect 30 340 64 345
rect 657 325 691 326
rect 542 -14 570 20
rect 605 -14 632 20
rect 1175 -14 1205 20
rect 1240 -14 1268 20
rect 1807 -14 1835 20
rect 1870 -14 1902 20
rect 2445 -14 2470 20
rect 2505 -14 2531 20
rect 2614 -14 2640 20
rect 2675 -14 2698 20
rect 3327 -14 3361 20
rect 3396 -14 3423 20
rect 4054 -14 4086 20
rect 4121 -14 4158 20
rect 4789 -14 4816 20
rect 4851 -14 4885 20
<< viali >>
rect 575 530 610 564
rect 1205 530 1240 564
rect 1840 530 1875 564
rect 2470 530 2505 564
rect 2640 530 2675 564
rect 3361 530 3396 564
rect 4091 530 4126 564
rect 4816 530 4851 564
rect 655 395 690 430
rect 25 305 60 340
rect 3261 310 3295 344
rect 3986 310 4020 344
rect 4716 310 4750 344
rect 5446 310 5480 344
rect 217 218 251 252
rect 345 218 379 252
rect 473 218 507 252
rect 852 218 886 252
rect 980 218 1014 252
rect 1108 218 1142 252
rect 1487 218 1521 252
rect 1615 218 1649 252
rect 1743 218 1777 252
rect 1925 225 1960 260
rect 2122 218 2156 252
rect 2250 218 2284 252
rect 2378 218 2412 252
rect 2779 218 2813 252
rect 2896 218 2930 252
rect 3504 218 3538 252
rect 3621 218 3655 252
rect 4234 218 4268 252
rect 4351 218 4385 252
rect 4964 218 4998 252
rect 5081 218 5115 252
rect 1295 120 1330 155
rect 570 -14 605 20
rect 1205 -14 1240 20
rect 1835 -14 1870 20
rect 2470 -14 2505 20
rect 2640 -14 2675 20
rect 3361 -14 3396 20
rect 4086 -14 4121 20
rect 4816 -14 4851 20
<< metal1 >>
rect 480 590 520 595
rect 541 564 631 595
rect 541 530 575 564
rect 610 530 631 564
rect 541 499 631 530
rect 1178 564 1270 595
rect 1178 530 1205 564
rect 1240 530 1270 564
rect 1178 499 1270 530
rect 1812 564 1902 595
rect 1812 530 1840 564
rect 1875 530 1902 564
rect 1812 499 1902 530
rect 2445 564 2529 595
rect 2445 530 2470 564
rect 2505 530 2529 564
rect 2445 499 2529 530
rect 2612 564 2701 595
rect 2612 530 2640 564
rect 2675 530 2701 564
rect 2612 499 2701 530
rect 3329 564 3423 595
rect 3329 530 3361 564
rect 3396 530 3423 564
rect 3329 499 3423 530
rect 4058 564 4153 595
rect 4058 530 4091 564
rect 4126 530 4153 564
rect 4058 499 4153 530
rect 4788 564 4885 595
rect 4788 530 4816 564
rect 4851 530 4885 564
rect 4788 499 4885 530
rect 635 445 715 455
rect 635 385 645 445
rect 705 385 715 445
rect 635 375 715 385
rect 3241 355 3321 365
rect 10 340 70 350
rect 10 305 25 340
rect 60 310 3180 340
rect 60 305 70 310
rect 10 290 70 305
rect 190 270 270 280
rect 190 210 200 270
rect 260 210 270 270
rect 190 200 270 210
rect 315 270 395 280
rect 315 210 325 270
rect 385 210 395 270
rect 315 200 395 210
rect 455 270 535 280
rect 980 275 1010 310
rect 455 210 465 270
rect 525 210 535 270
rect 455 200 535 210
rect 825 265 905 275
rect 825 205 835 265
rect 895 205 905 265
rect 825 195 905 205
rect 955 265 1035 275
rect 955 205 965 265
rect 1025 205 1035 265
rect 955 195 1035 205
rect 1085 265 1165 275
rect 1085 205 1095 265
rect 1155 205 1165 265
rect 1085 195 1165 205
rect 1460 265 1540 275
rect 1460 205 1470 265
rect 1530 205 1540 265
rect 1460 195 1540 205
rect 1585 265 1665 275
rect 1585 205 1595 265
rect 1655 205 1665 265
rect 1585 195 1665 205
rect 1725 265 1805 275
rect 1725 205 1735 265
rect 1795 205 1805 265
rect 1725 195 1805 205
rect 1905 265 1985 275
rect 1905 205 1915 265
rect 1975 205 1985 265
rect 1905 195 1985 205
rect 2095 265 2175 275
rect 2095 205 2105 265
rect 2165 205 2175 265
rect 2095 195 2175 205
rect 2230 265 2310 275
rect 2230 205 2240 265
rect 2300 205 2310 265
rect 2230 195 2310 205
rect 2360 265 2440 275
rect 2360 205 2370 265
rect 2430 205 2440 265
rect 2360 195 2440 205
rect 2756 260 2836 270
rect 2756 200 2766 260
rect 2826 200 2836 260
rect 1280 155 1340 165
rect 2250 155 2280 195
rect 2756 190 2836 200
rect 2876 265 2956 275
rect 2876 205 2886 265
rect 2946 205 2956 265
rect 3150 250 3180 310
rect 3241 295 3251 355
rect 3311 295 3321 355
rect 3241 285 3321 295
rect 3966 350 4046 360
rect 3966 295 3976 350
rect 4036 295 4046 350
rect 3966 285 4046 295
rect 4696 355 4776 365
rect 4696 295 4706 355
rect 4766 295 4776 355
rect 4696 285 4776 295
rect 5426 355 5506 365
rect 5426 300 5436 355
rect 5496 300 5506 355
rect 5426 290 5506 300
rect 3481 270 3561 280
rect 3481 250 3491 270
rect 3150 220 3491 250
rect 2876 195 2956 205
rect 3481 210 3491 220
rect 3551 210 3561 270
rect 4211 265 4291 275
rect 3481 200 3561 210
rect 3596 255 3676 265
rect 3596 195 3606 255
rect 3666 195 3676 255
rect 4211 205 4221 265
rect 4281 205 4291 265
rect 4211 195 4291 205
rect 4326 265 4406 275
rect 4326 205 4336 265
rect 4396 205 4406 265
rect 4326 195 4406 205
rect 4941 265 5021 275
rect 4941 205 4951 265
rect 5011 205 5021 265
rect 4941 195 5021 205
rect 5056 265 5136 275
rect 5056 205 5066 265
rect 5126 205 5136 265
rect 5056 195 5136 205
rect 3596 185 3676 195
rect 4965 155 4995 195
rect 1280 120 1295 155
rect 1330 125 4995 155
rect 1330 120 1340 125
rect 1280 105 1340 120
rect 539 20 636 51
rect 539 -14 570 20
rect 605 -14 636 20
rect 539 -45 636 -14
rect 1167 20 1269 51
rect 1167 -14 1205 20
rect 1240 -14 1269 20
rect 1167 -45 1269 -14
rect 1813 20 1901 51
rect 1813 -14 1835 20
rect 1870 -14 1901 20
rect 1813 -45 1901 -14
rect 2438 20 2534 51
rect 2438 -14 2470 20
rect 2505 -14 2534 20
rect 2438 -45 2534 -14
rect 2608 20 2698 51
rect 2608 -14 2640 20
rect 2675 -14 2698 20
rect 2608 -45 2698 -14
rect 3334 20 3424 51
rect 3334 -14 3361 20
rect 3396 -14 3424 20
rect 3334 -45 3424 -14
rect 4058 20 4154 51
rect 4058 -14 4086 20
rect 4121 -14 4154 20
rect 4058 -45 4154 -14
rect 4788 20 4885 51
rect 4788 -14 4816 20
rect 4851 -14 4885 20
rect 4788 -45 4885 -14
rect 450 -85 530 -75
rect 450 -145 460 -85
rect 520 -100 530 -85
rect 2875 -85 2955 -75
rect 2875 -100 2885 -85
rect 520 -130 2885 -100
rect 520 -145 530 -130
rect 450 -155 530 -145
rect 2875 -145 2885 -130
rect 2945 -145 2955 -85
rect 2875 -155 2955 -145
rect 1085 -170 1165 -160
rect 1085 -230 1095 -170
rect 1155 -185 1165 -170
rect 3595 -170 3675 -160
rect 3595 -185 3605 -170
rect 1155 -215 3605 -185
rect 1155 -230 1165 -215
rect 1085 -240 1165 -230
rect 3595 -230 3605 -215
rect 3665 -230 3675 -170
rect 3595 -240 3675 -230
rect 1720 -255 1800 -245
rect 1720 -315 1730 -255
rect 1790 -270 1800 -255
rect 4330 -255 4410 -245
rect 4330 -270 4340 -255
rect 1790 -300 4340 -270
rect 1790 -315 1800 -300
rect 1720 -325 1800 -315
rect 4330 -315 4340 -300
rect 4400 -315 4410 -255
rect 4330 -325 4410 -315
rect 2355 -340 2435 -330
rect 2355 -400 2365 -340
rect 2425 -355 2435 -340
rect 5060 -340 5140 -330
rect 5060 -355 5070 -340
rect 2425 -385 5070 -355
rect 2425 -400 2435 -385
rect 2355 -410 2435 -400
rect 5060 -400 5070 -385
rect 5130 -400 5140 -340
rect 5060 -410 5140 -400
rect 325 -425 410 -415
rect 325 -485 335 -425
rect 400 -440 410 -425
rect 2755 -425 2835 -415
rect 2755 -440 2765 -425
rect 400 -470 2765 -440
rect 400 -485 410 -470
rect 325 -495 410 -485
rect 2755 -485 2765 -470
rect 2825 -485 2835 -425
rect 2755 -495 2835 -485
rect 630 -510 710 -500
rect 630 -570 640 -510
rect 700 -525 710 -510
rect 1590 -510 1670 -500
rect 1590 -525 1600 -510
rect 700 -555 1600 -525
rect 700 -570 710 -555
rect 630 -580 710 -570
rect 1590 -570 1600 -555
rect 1660 -525 1670 -510
rect 4210 -510 4290 -500
rect 4210 -525 4220 -510
rect 1660 -555 4220 -525
rect 1660 -570 1670 -555
rect 1590 -580 1670 -570
rect 4210 -570 4220 -555
rect 4280 -570 4290 -510
rect 4210 -580 4290 -570
<< via1 >>
rect 645 430 705 445
rect 645 395 655 430
rect 655 395 690 430
rect 690 395 705 430
rect 645 385 705 395
rect 200 252 260 270
rect 200 218 217 252
rect 217 218 251 252
rect 251 218 260 252
rect 200 210 260 218
rect 325 252 385 270
rect 325 218 345 252
rect 345 218 379 252
rect 379 218 385 252
rect 325 210 385 218
rect 465 252 525 270
rect 465 218 473 252
rect 473 218 507 252
rect 507 218 525 252
rect 465 210 525 218
rect 835 252 895 265
rect 835 218 852 252
rect 852 218 886 252
rect 886 218 895 252
rect 835 205 895 218
rect 965 252 1025 265
rect 965 218 980 252
rect 980 218 1014 252
rect 1014 218 1025 252
rect 965 205 1025 218
rect 1095 252 1155 265
rect 1095 218 1108 252
rect 1108 218 1142 252
rect 1142 218 1155 252
rect 1095 205 1155 218
rect 1470 252 1530 265
rect 1470 218 1487 252
rect 1487 218 1521 252
rect 1521 218 1530 252
rect 1470 205 1530 218
rect 1595 252 1655 265
rect 1595 218 1615 252
rect 1615 218 1649 252
rect 1649 218 1655 252
rect 1595 205 1655 218
rect 1735 252 1795 265
rect 1735 218 1743 252
rect 1743 218 1777 252
rect 1777 218 1795 252
rect 1735 205 1795 218
rect 1915 260 1975 265
rect 1915 225 1925 260
rect 1925 225 1960 260
rect 1960 225 1975 260
rect 1915 205 1975 225
rect 2105 252 2165 265
rect 2105 218 2122 252
rect 2122 218 2156 252
rect 2156 218 2165 252
rect 2105 205 2165 218
rect 2240 252 2300 265
rect 2240 218 2250 252
rect 2250 218 2284 252
rect 2284 218 2300 252
rect 2240 205 2300 218
rect 2370 252 2430 265
rect 2370 218 2378 252
rect 2378 218 2412 252
rect 2412 218 2430 252
rect 2370 205 2430 218
rect 2766 252 2826 260
rect 2766 218 2779 252
rect 2779 218 2813 252
rect 2813 218 2826 252
rect 2766 200 2826 218
rect 2886 252 2946 265
rect 2886 218 2896 252
rect 2896 218 2930 252
rect 2930 218 2946 252
rect 2886 205 2946 218
rect 3251 344 3311 355
rect 3251 310 3261 344
rect 3261 310 3295 344
rect 3295 310 3311 344
rect 3251 295 3311 310
rect 3976 344 4036 350
rect 3976 310 3986 344
rect 3986 310 4020 344
rect 4020 310 4036 344
rect 3976 295 4036 310
rect 4706 344 4766 355
rect 4706 310 4716 344
rect 4716 310 4750 344
rect 4750 310 4766 344
rect 4706 295 4766 310
rect 5436 344 5496 355
rect 5436 310 5446 344
rect 5446 310 5480 344
rect 5480 310 5496 344
rect 5436 300 5496 310
rect 3491 252 3551 270
rect 3491 218 3504 252
rect 3504 218 3538 252
rect 3538 218 3551 252
rect 3491 210 3551 218
rect 3606 252 3666 255
rect 3606 218 3621 252
rect 3621 218 3655 252
rect 3655 218 3666 252
rect 3606 195 3666 218
rect 4221 252 4281 265
rect 4221 218 4234 252
rect 4234 218 4268 252
rect 4268 218 4281 252
rect 4221 205 4281 218
rect 4336 252 4396 265
rect 4336 218 4351 252
rect 4351 218 4385 252
rect 4385 218 4396 252
rect 4336 205 4396 218
rect 4951 252 5011 265
rect 4951 218 4964 252
rect 4964 218 4998 252
rect 4998 218 5011 252
rect 4951 205 5011 218
rect 5066 252 5126 265
rect 5066 218 5081 252
rect 5081 218 5115 252
rect 5115 218 5126 252
rect 5066 205 5126 218
rect 460 -145 520 -85
rect 2885 -145 2945 -85
rect 1095 -230 1155 -170
rect 3605 -230 3665 -170
rect 1730 -315 1790 -255
rect 4340 -315 4400 -255
rect 2365 -400 2425 -340
rect 5070 -400 5130 -340
rect 335 -485 400 -425
rect 2765 -485 2825 -425
rect 640 -570 700 -510
rect 1600 -570 1660 -510
rect 4220 -570 4280 -510
<< metal2 >>
rect 635 445 715 455
rect 635 385 645 445
rect 705 385 715 445
rect 635 375 715 385
rect 190 270 270 280
rect 190 210 200 270
rect 260 210 270 270
rect 190 200 270 210
rect 315 270 395 280
rect 315 210 325 270
rect 385 210 395 270
rect 315 200 395 210
rect 455 270 535 280
rect 455 210 465 270
rect 525 210 535 270
rect 455 200 535 210
rect 350 -415 380 200
rect 475 -75 505 200
rect 450 -85 530 -75
rect 450 -145 460 -85
rect 520 -145 530 -85
rect 450 -155 530 -145
rect 325 -425 410 -415
rect 325 -485 335 -425
rect 400 -485 410 -425
rect 325 -495 410 -485
rect 655 -500 685 375
rect 3241 355 3321 365
rect 3241 295 3251 355
rect 3311 295 3321 355
rect 3241 285 3321 295
rect 3966 350 4046 360
rect 3966 295 3976 350
rect 4036 295 4046 350
rect 3966 285 4046 295
rect 4696 355 4776 365
rect 4696 295 4706 355
rect 4766 295 4776 355
rect 4696 285 4776 295
rect 5426 355 5506 365
rect 5426 300 5436 355
rect 5496 300 5506 355
rect 5426 290 5506 300
rect 825 265 905 275
rect 825 205 835 265
rect 895 205 905 265
rect 825 195 905 205
rect 955 265 1035 275
rect 955 205 965 265
rect 1025 205 1035 265
rect 955 195 1035 205
rect 1085 265 1165 275
rect 1085 205 1095 265
rect 1155 205 1165 265
rect 1085 195 1165 205
rect 1460 265 1540 275
rect 1460 205 1470 265
rect 1530 205 1540 265
rect 1460 195 1540 205
rect 1585 265 1665 275
rect 1585 205 1595 265
rect 1655 205 1665 265
rect 1585 195 1665 205
rect 1725 265 1805 275
rect 1725 205 1735 265
rect 1795 205 1805 265
rect 1110 -160 1140 195
rect 1085 -170 1165 -160
rect 1085 -230 1095 -170
rect 1155 -230 1165 -170
rect 1085 -240 1165 -230
rect 1615 -500 1645 195
rect 1725 194 1805 205
rect 1905 265 1985 275
rect 1905 205 1915 265
rect 1975 205 1985 265
rect 1905 195 1985 205
rect 2095 265 2175 275
rect 2095 205 2105 265
rect 2165 205 2175 265
rect 2095 195 2175 205
rect 2230 265 2310 275
rect 2230 205 2240 265
rect 2300 205 2310 265
rect 2230 195 2310 205
rect 2360 265 2440 275
rect 2360 205 2370 265
rect 2430 205 2440 265
rect 2360 195 2440 205
rect 2756 260 2836 270
rect 2756 200 2766 260
rect 2826 200 2836 260
rect 1745 -245 1775 194
rect 1720 -255 1800 -245
rect 1720 -315 1730 -255
rect 1790 -315 1800 -255
rect 1720 -325 1800 -315
rect 2380 -330 2410 195
rect 2756 190 2836 200
rect 2876 265 2956 275
rect 2876 205 2886 265
rect 2946 205 2956 265
rect 2876 195 2956 205
rect 3481 270 3561 280
rect 3481 210 3491 270
rect 3551 210 3561 270
rect 4211 265 4291 275
rect 3481 200 3561 210
rect 3596 255 3676 265
rect 3596 195 3606 255
rect 3666 195 3676 255
rect 4211 205 4221 265
rect 4281 205 4291 265
rect 4211 195 4291 205
rect 4326 265 4406 275
rect 4326 205 4336 265
rect 4396 205 4406 265
rect 4326 195 4406 205
rect 4941 265 5021 275
rect 4941 205 4951 265
rect 5011 205 5021 265
rect 4941 195 5021 205
rect 5056 265 5136 275
rect 5056 205 5066 265
rect 5126 205 5136 265
rect 5056 195 5136 205
rect 2355 -340 2435 -330
rect 2355 -400 2365 -340
rect 2425 -400 2435 -340
rect 2355 -410 2435 -400
rect 2780 -415 2810 190
rect 2900 -75 2930 195
rect 3596 185 3676 195
rect 2875 -85 2955 -75
rect 2875 -145 2885 -85
rect 2945 -145 2955 -85
rect 2875 -155 2955 -145
rect 3620 -160 3650 185
rect 3595 -170 3675 -160
rect 3595 -230 3605 -170
rect 3665 -230 3675 -170
rect 3595 -240 3675 -230
rect 2755 -425 2835 -415
rect 2755 -485 2765 -425
rect 2825 -485 2835 -425
rect 2755 -495 2835 -485
rect 4235 -500 4265 195
rect 4355 -245 4385 195
rect 4330 -255 4410 -245
rect 4330 -315 4340 -255
rect 4400 -315 4410 -255
rect 4330 -325 4410 -315
rect 5085 -330 5115 195
rect 5060 -340 5140 -330
rect 5060 -400 5070 -340
rect 5130 -400 5140 -340
rect 5060 -410 5140 -400
rect 630 -510 710 -500
rect 630 -570 640 -510
rect 700 -570 710 -510
rect 630 -580 710 -570
rect 1590 -510 1670 -500
rect 1590 -570 1600 -510
rect 1660 -570 1670 -510
rect 1590 -580 1670 -570
rect 4210 -510 4290 -500
rect 4210 -570 4220 -510
rect 4280 -570 4290 -510
rect 4210 -580 4290 -570
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_0
timestamp 1691611044
transform 1 0 -7 0 1 3
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_1
timestamp 1691611044
transform 1 0 628 0 1 3
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_2
timestamp 1691611044
transform 1 0 1263 0 1 3
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  sky130_fd_sc_hd__a21o_1_3
timestamp 1691611044
transform 1 0 1898 0 1 3
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  sky130_fd_sc_hd__tapvpwrvgnd_1_0
timestamp 1691611044
transform 1 0 2526 0 1 3
box -38 -48 130 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_0
timestamp 1691611044
transform 1 0 2694 0 1 3
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_1
timestamp 1691611044
transform 1 0 3419 0 1 3
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_2
timestamp 1691611044
transform 1 0 4149 0 1 3
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  sky130_fd_sc_hd__xor2_1_3
timestamp 1691611044
transform 1 0 4879 0 1 3
box -38 -48 682 592
<< labels >>
flabel via1 490 240 490 240 1 FreeSans 128 0 0 0 P1
port 2 n
flabel via1 360 240 360 240 1 FreeSans 160 0 0 0 CI
port 1 n
flabel via1 1125 235 1125 235 1 FreeSans 240 0 0 0 P2
port 4 n
flabel via1 234 240 234 240 1 FreeSans 128 0 0 0 G1
port 3 n
flabel via1 870 240 870 240 1 FreeSans 160 0 0 0 G2
port 5 n
flabel via1 1760 245 1760 245 1 FreeSans 128 0 0 0 P3
port 6 n
flabel via1 1500 245 1500 245 1 FreeSans 128 0 0 0 G3
port 7 n
flabel via1 2395 241 2395 241 1 FreeSans 128 0 0 0 P4
port 8 n
flabel via1 2138 240 2138 240 1 FreeSans 128 0 0 0 G4
port 9 n
flabel via1 1935 240 1935 240 1 FreeSans 160 0 0 0 CO
port 14 n
flabel via1 4001 335 4001 335 1 FreeSans 128 0 0 0 S2
port 11 n
flabel via1 4731 335 4731 335 1 FreeSans 160 0 0 0 S3
port 12 n
flabel via1 5461 335 5461 335 1 FreeSans 160 0 0 0 S4
port 13 n
flabel via1 3276 335 3276 335 1 FreeSans 128 0 0 0 S1
port 10 n
flabel nwell s 2565 350 2565 350 1 FreeSans 240 0 0 0 VPB
port 17 n
flabel pwell s 2565 120 2565 120 1 FreeSans 240 0 0 0 VNB
port 18 n
flabel metal1 s 555 35 555 35 1 FreeSans 160 0 0 0 GND
port 16 n
flabel viali s 595 550 595 550 1 FreeSans 160 0 0 0 VDD
port 15 n
<< end >>
